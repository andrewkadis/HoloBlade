// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Fri Aug 28 18:30:53 2020
//
// Verilog Description of module top
//

module top (ICE_SYSCLK, DCD, DSR, DTR, CTS, RST, UART_RX, UART_TX, 
            SEN, SCK, SOUT, SDAT, UPDATE, RESET, SLM_CLK, INVERT, 
            SYNC, VALID, DATA31, DATA0, DATA30, DATA29, DATA1, 
            DATA28, DATA27, DATA2, DATA26, DATA25, DATA3, DATA24, 
            DATA23, DATA4, DATA22, DATA21, DATA5, DATA20, DATA19, 
            DATA6, DATA18, DATA17, DATA7, DATA16, DATA15, DATA8, 
            DATA14, DATA13, DATA12, DATA11, DATA9, DATA10, FT_OE, 
            FT_RD, FT_WR, FT_SIWU, FR_RXF, FT_TXE, FIFO_BE3, FIFO_BE2, 
            FIFO_BE1, FIFO_BE0, FIFO_D31, FIFO_D30, FIFO_D29, FIFO_D28, 
            FIFO_D27, FIFO_CLK, FIFO_D26, FIFO_D25, FIFO_D24, FIFO_D23, 
            FIFO_D22, FIFO_D21, FIFO_D20, FIFO_D19, FIFO_D18, FIFO_D17, 
            FIFO_D16, FIFO_D15, FIFO_D14, FIFO_D13, FIFO_D12, FIFO_D11, 
            FIFO_D10, FIFO_D9, FIFO_D8, FIFO_D7, FIFO_D6, FIFO_D5, 
            FIFO_D4, FIFO_D3, FIFO_D2, FIFO_D1, FIFO_D0, DEBUG_0, 
            DEBUG_1, DEBUG_2, DEBUG_3, DEBUG_5, DEBUG_6, DEBUG_8, 
            DEBUG_9, ICE_CLK, ICE_CDONE, ICE_CREST) /* synthesis syn_module_defined=1 */ ;   // src/top.v(5[8:11])
    input ICE_SYSCLK;   // src/top.v(8[11:21])
    output DCD;   // src/top.v(11[12:15])
    output DSR;   // src/top.v(12[12:15])
    output DTR;   // src/top.v(13[12:15])
    output CTS;   // src/top.v(14[12:15])
    output RST;   // src/top.v(15[12:15])
    input UART_RX;   // src/top.v(16[12:19])
    output UART_TX;   // src/top.v(17[12:19])
    output SEN;   // src/top.v(20[12:15])
    output SCK;   // src/top.v(21[12:15])
    input SOUT;   // src/top.v(22[12:16])
    output SDAT;   // src/top.v(23[12:16])
    output UPDATE;   // src/top.v(27[12:18])
    output RESET;   // src/top.v(28[12:17])
    output SLM_CLK;   // src/top.v(29[12:19])
    output INVERT;   // src/top.v(30[12:18])
    output SYNC;   // src/top.v(31[12:16])
    output VALID;   // src/top.v(32[12:17])
    output DATA31;   // src/top.v(34[12:18])
    output DATA0;   // src/top.v(35[12:17])
    output DATA30;   // src/top.v(36[12:18])
    output DATA29;   // src/top.v(37[12:18])
    output DATA1;   // src/top.v(38[12:17])
    output DATA28;   // src/top.v(39[12:18])
    output DATA27;   // src/top.v(40[12:18])
    output DATA2;   // src/top.v(41[12:17])
    output DATA26;   // src/top.v(42[12:18])
    output DATA25;   // src/top.v(43[12:18])
    output DATA3;   // src/top.v(44[12:17])
    output DATA24;   // src/top.v(45[12:18])
    output DATA23;   // src/top.v(46[12:18])
    output DATA4;   // src/top.v(47[12:17])
    output DATA22;   // src/top.v(48[12:18])
    output DATA21;   // src/top.v(49[12:18])
    output DATA5;   // src/top.v(50[12:17])
    output DATA20;   // src/top.v(51[12:18])
    output DATA19;   // src/top.v(52[12:18])
    output DATA6;   // src/top.v(53[12:17])
    output DATA18;   // src/top.v(54[12:18])
    output DATA17;   // src/top.v(55[12:18])
    output DATA7;   // src/top.v(56[12:17])
    output DATA16;   // src/top.v(57[12:18])
    output DATA15;   // src/top.v(58[12:18])
    output DATA8;   // src/top.v(59[12:17])
    output DATA14;   // src/top.v(60[12:18])
    output DATA13;   // src/top.v(61[12:18])
    output DATA12;   // src/top.v(62[12:18])
    output DATA11;   // src/top.v(63[12:18])
    output DATA9;   // src/top.v(64[12:17])
    output DATA10;   // src/top.v(65[12:18])
    output FT_OE;   // src/top.v(69[12:17])
    output FT_RD;   // src/top.v(70[12:17])
    output FT_WR;   // src/top.v(71[12:17])
    output FT_SIWU;   // src/top.v(72[12:19])
    input FR_RXF;   // src/top.v(73[12:18])
    input FT_TXE;   // src/top.v(74[12:18])
    input FIFO_BE3;   // src/top.v(75[12:20])
    input FIFO_BE2;   // src/top.v(76[12:20])
    input FIFO_BE1;   // src/top.v(77[12:20])
    input FIFO_BE0;   // src/top.v(78[12:20])
    input FIFO_D31;   // src/top.v(79[12:20])
    input FIFO_D30;   // src/top.v(80[12:20])
    input FIFO_D29;   // src/top.v(81[12:20])
    input FIFO_D28;   // src/top.v(82[12:20])
    input FIFO_D27;   // src/top.v(83[12:20])
    input FIFO_CLK;   // src/top.v(84[12:20])
    input FIFO_D26;   // src/top.v(85[12:20])
    input FIFO_D25;   // src/top.v(86[12:20])
    input FIFO_D24;   // src/top.v(87[12:20])
    input FIFO_D23;   // src/top.v(88[12:20])
    input FIFO_D22;   // src/top.v(89[12:20])
    input FIFO_D21;   // src/top.v(90[12:20])
    input FIFO_D20;   // src/top.v(91[12:20])
    input FIFO_D19;   // src/top.v(92[12:20])
    input FIFO_D18;   // src/top.v(93[12:20])
    input FIFO_D17;   // src/top.v(94[12:20])
    input FIFO_D16;   // src/top.v(95[12:20])
    input FIFO_D15;   // src/top.v(97[11:19])
    input FIFO_D14;   // src/top.v(98[11:19])
    input FIFO_D13;   // src/top.v(99[11:19])
    input FIFO_D12;   // src/top.v(100[11:19])
    input FIFO_D11;   // src/top.v(101[11:19])
    input FIFO_D10;   // src/top.v(102[11:19])
    input FIFO_D9;   // src/top.v(103[11:18])
    input FIFO_D8;   // src/top.v(104[11:18])
    input FIFO_D7;   // src/top.v(105[11:18])
    input FIFO_D6;   // src/top.v(106[11:18])
    input FIFO_D5;   // src/top.v(107[11:18])
    input FIFO_D4;   // src/top.v(108[11:18])
    input FIFO_D3;   // src/top.v(109[11:18])
    input FIFO_D2;   // src/top.v(110[11:18])
    input FIFO_D1;   // src/top.v(111[11:18])
    input FIFO_D0;   // src/top.v(112[11:18])
    output DEBUG_0;   // src/top.v(115[12:19])
    output DEBUG_1;   // src/top.v(116[12:19])
    output DEBUG_2;   // src/top.v(117[12:19])
    output DEBUG_3;   // src/top.v(118[12:19])
    output DEBUG_5;   // src/top.v(119[12:19])
    output DEBUG_6;   // src/top.v(120[12:19])
    output DEBUG_8;   // src/top.v(121[12:19])
    output DEBUG_9;   // src/top.v(122[12:19])
    output ICE_CLK;   // src/top.v(125[12:19])
    output ICE_CDONE;   // src/top.v(126[12:21])
    output ICE_CREST;   // src/top.v(127[12:21])
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    
    wire GND_net, VCC_net, ICE_SYSCLK_c, UART_RX_c, UART_TX_c, SEN_c_1, 
        SCK_c_0, SOUT_c, SDAT_c_15, UPDATE_c_2, RESET_c, INVERT_c_3, 
        SYNC_c, DEBUG_9_c, DATA15_c, DEBUG_6_c, DATA14_c, DATA13_c, 
        DATA17_c, DATA12_c, DATA11_c, DATA18_c, DATA10_c, DATA9_c, 
        DATA19_c, DATA8_c, DATA7_c, DATA20_c, DATA6_c, DATA5_c, 
        FT_OE_c, DEBUG_2_c, DEBUG_1_c_c, FIFO_D15_c_15, FIFO_D14_c_14, 
        FIFO_D13_c_13, FIFO_D12_c_12, FIFO_D11_c_11, FIFO_D10_c_10, 
        FIFO_D9_c_9, FIFO_D8_c_8, FIFO_D7_c_7, FIFO_D6_c_6, FIFO_D5_c_5, 
        FIFO_D4_c_4, FIFO_D3_c_3, FIFO_D2_c_2, FIFO_D1_c_1, DEBUG_8_c_0_c, 
        DEBUG_0_c_24, DEBUG_3_c, DEBUG_5_c, debug_led3, reset_all_w;
    wire [3:0]reset_clk_counter;   // src/top.v(242[10:27])
    
    wire reset_per_frame, buffer_switch_done, dc32_fifo_almost_full, \REG.mem_13_13 , 
        \REG.mem_13_12 , \REG.mem_13_11 , \REG.mem_13_10 , \REG.mem_13_9 , 
        \REG.mem_13_8 , \REG.mem_13_7 , \REG.mem_13_6 , \REG.mem_11_15 , 
        \REG.mem_11_14 , \REG.mem_11_13 , \REG.mem_11_12 , \REG.mem_11_11 , 
        \REG.mem_11_10 , \REG.mem_11_9 ;
    wire [31:0]dc32_fifo_data_in;   // src/top.v(510[13:30])
    
    wire dc32_fifo_almost_empty, get_next_word, \REG.mem_9_14 , \REG.mem_9_13 , 
        \REG.mem_9_12 , \REG.mem_9_11 , \REG.mem_9_10 , \REG.mem_9_9 , 
        \REG.mem_9_8 , \REG.mem_9_7 , \REG.mem_9_6 , \REG.mem_9_5 , 
        \REG.mem_9_4 , \REG.mem_9_3 , \REG.mem_9_2 , \REG.mem_9_1 , 
        \REG.mem_9_0 ;
    wire [31:0]fifo_data_out;   // src/top.v(545[12:25])
    wire [7:0]pc_data_rx;   // src/top.v(685[11:21])
    
    wire \REG.mem_15_15 , tx_uart_active_flag, spi_start_transfer_r, multi_byte_spi_trans_flag_r;
    wire [7:0]tx_addr_byte;   // src/top.v(807[11:23])
    wire [7:0]tx_data_byte;   // src/top.v(809[11:23])
    wire [7:0]rx_buf_byte;   // src/top.v(816[11:22])
    
    wire is_tx_fifo_full_flag, fifo_write_cmd, spi_rx_byte_ready, fifo_read_cmd, 
        is_fifo_empty_flag;
    wire [31:0]fifo_temp_output;   // src/top.v(906[12:28])
    
    wire even_byte_flag, uart_rx_complete_rising_edge, uart_rx_complete_prev, 
        \REG.mem_15_14 , reset_all_w_N_61, \REG.mem_11_8 , \REG.mem_11_7 , 
        start_tx_N_64, pll_clk_unbuf, n7386;
    wire [3:0]state;   // src/timing_controller.v(51[11:16])
    
    wire n771, multi_byte_spi_trans_flag_r_N_72, \REG.mem_8_15 , \REG.mem_18_15 , 
        \REG.mem_18_14 , \REG.mem_18_13 , \REG.mem_18_12 , \REG.mem_18_11 , 
        \REG.mem_18_10 , \REG.mem_18_9 , \REG.mem_18_8 , \REG.mem_18_7 , 
        \REG.mem_18_6 , \REG.mem_18_5 , \REG.mem_18_4 , \REG.mem_18_3 , 
        \REG.mem_18_2 , \REG.mem_18_1 , \REG.mem_18_0 , n4253, \REG.mem_16_15 , 
        \REG.mem_16_14 , \REG.mem_16_13 , \REG.mem_16_12 , \REG.mem_16_11 , 
        \REG.mem_16_10 , \REG.mem_16_9 , \REG.mem_16_8 , \REG.mem_16_7 , 
        \REG.mem_16_6 , \REG.mem_16_5 , \REG.mem_16_4 , \REG.mem_16_3 , 
        \REG.mem_16_2 , \REG.mem_8_14 , \REG.mem_8_13 , \REG.mem_8_12 , 
        \REG.mem_8_11 , \REG.mem_8_10 , \REG.mem_8_9 , \REG.mem_8_8 , 
        \REG.mem_8_7 , \REG.mem_8_6 , \REG.mem_8_5 , \REG.mem_8_4 , 
        \REG.mem_8_3 , \REG.mem_8_2 , \REG.mem_8_1 , \REG.mem_8_0 , 
        \REG.mem_7_15 , \REG.mem_15_13 , reset_per_frame_latched, \REG.mem_11_6 , 
        buffer_switch_done_latched, \REG.mem_11_5 , \REG.mem_11_4 , \REG.mem_11_3 , 
        \REG.mem_11_2 , \REG.mem_11_1 , \REG.mem_11_0 , n2352, \REG.mem_16_1 , 
        \REG.mem_16_0 , n2034, n2086, n4942, n4939, \REG.mem_12_2 , 
        \REG.mem_12_3 , write_to_dc32_fifo_latched_N_425, FT_OE_N_420, 
        \REG.mem_10_15 , \REG.mem_10_14 , \REG.mem_10_13 , n4937, \REG.mem_10_12 , 
        n4936, \REG.mem_10_11 , \REG.mem_10_10 , \REG.mem_10_9 , \REG.mem_10_8 , 
        \REG.mem_10_7 , \REG.mem_10_6 , \REG.mem_14_11 , \REG.mem_14_12 , 
        \REG.mem_14_13 , \REG.mem_14_14 , \REG.mem_14_15 , \REG.mem_10_5 , 
        \REG.mem_10_4 , \REG.mem_10_3 , \REG.mem_10_2 , \REG.mem_10_1 , 
        \REG.mem_10_0 , \REG.mem_15_12 , \REG.mem_15_11 , \REG.mem_15_10 , 
        \REG.mem_15_9 , n4923, n4922, n4919, \REG.mem_9_15 , \REG.mem_3_0 , 
        \REG.mem_7_14 , \REG.mem_7_13 , \REG.mem_7_12 , \REG.mem_7_11 , 
        \REG.mem_13_5 , \REG.mem_15_8 , \REG.mem_15_7 , \REG.mem_15_6 , 
        \REG.mem_13_0 , n4916, n4911, n4910, n4909, \REG.mem_15_5 , 
        n4907, n4904, n4903, n4901, n4899, n4898, n4897, \REG.mem_7_10 , 
        \REG.mem_7_9 , \REG.mem_7_8 , \REG.mem_7_7 , \REG.mem_7_6 , 
        \REG.mem_7_5 , \REG.mem_7_4 , \REG.mem_7_3 , bluejay_data_out_31__N_736, 
        bluejay_data_out_31__N_737, n575, r_Rx_Data;
    wire [2:0]r_SM_Main;   // src/uart_rx.v(36[17:26])
    
    wire n1879, \REG.mem_12_1 , \REG.mem_12_0 , \REG.mem_15_4 , \REG.mem_14_10 , 
        \REG.mem_14_8 , \REG.mem_14_7 , \REG.mem_15_3 ;
    wire [2:0]r_SM_Main_2__N_765;
    
    wire n4661;
    wire [2:0]r_SM_Main_adj_95;   // src/uart_tx.v(31[16:25])
    wire [7:0]r_Tx_Data;   // src/uart_tx.v(34[16:25])
    
    wire n10277;
    wire [2:0]r_SM_Main_2__N_844;
    wire [2:0]r_SM_Main_2__N_841;
    
    wire \REG.mem_15_2 , \REG.mem_14_6 , \REG.mem_14_5 , \REG.mem_15_1 , 
        n10428, \REG.mem_14_9 ;
    wire [15:0]tx_shift_reg;   // src/spi.v(70[12:24])
    wire [15:0]rx_shift_reg;   // src/spi.v(72[12:24])
    
    wire \REG.mem_15_0 , n4245, n4890, n4889, n571, n4888, n4887, 
        n4883, n4882, \REG.mem_7_2 , \REG.mem_7_1 , \REG.mem_7_0 , 
        \REG.mem_14_2 , \REG.mem_14_1 , \REG.mem_14_3 , \REG.mem_14_4 , 
        \REG.mem_6_15 , \REG.mem_6_14 , \REG.mem_6_13 , \REG.mem_6_12 , 
        \REG.mem_6_11 , \REG.mem_6_10 , \REG.mem_6_9 , \REG.mem_6_8 , 
        \REG.mem_6_7 , \REG.mem_6_6 , \REG.mem_6_5 , \REG.mem_6_4 , 
        \REG.mem_6_3 , \REG.mem_6_2 , \REG.mem_6_1 , \REG.mem_6_0 , 
        \REG.mem_13_1 , \REG.mem_13_15 , \REG.mem_13_2 , \REG.mem_13_3 ;
    wire [6:0]wr_addr_nxt_c;   // src/fifo_dc_32_lut_gen.v(198[29:42])
    wire [6:0]rp_sync1_r;   // src/fifo_dc_32_lut_gen.v(201[37:47])
    wire [6:0]wr_grey_sync_r;   // src/fifo_dc_32_lut_gen.v(204[37:51])
    wire [6:0]rd_addr_r;   // src/fifo_dc_32_lut_gen.v(217[29:38])
    
    wire \REG.mem_14_0 ;
    wire [6:0]rd_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(221[30:42])
    wire [6:0]wp_sync1_r;   // src/fifo_dc_32_lut_gen.v(222[37:47])
    wire [6:0]rd_grey_sync_r;   // src/fifo_dc_32_lut_gen.v(225[37:51])
    wire [6:0]rd_sig_diff0_w;   // src/fifo_dc_32_lut_gen.v(233[30:44])
    
    wire rd_fifo_en_w, \aempty_flag_impl.ae_flag_nxt_w , t_rd_fifo_en_w;
    wire [31:0]\REG.out_raw ;   // src/fifo_dc_32_lut_gen.v(879[47:54])
    wire [6:0]rd_addr_nxt_c_6__N_498;
    
    wire n4, n7590, \REG.mem_5_15 , \REG.mem_5_14 , \REG.mem_5_13 , 
        \REG.mem_5_12 , \REG.mem_5_11 , \REG.mem_5_10 , \REG.mem_5_9 , 
        \REG.mem_5_8 , \REG.mem_5_7 , \REG.mem_5_6 , \REG.mem_5_5 , 
        \REG.mem_5_4 , \REG.mem_5_3 , \REG.mem_5_2 , \REG.mem_5_1 , 
        \REG.mem_5_0 , n8, n4878, n7568, n4877, \REG.mem_4_15 , 
        \REG.mem_4_14 , \REG.mem_4_13 , \REG.mem_4_12 , \REG.mem_4_11 , 
        \REG.mem_4_10 , \REG.mem_4_9 , \REG.mem_4_8 , \REG.mem_4_7 , 
        \REG.mem_4_6 , \REG.mem_4_5 , \REG.mem_4_4 , \REG.mem_4_3 , 
        \REG.mem_4_2 , \REG.mem_4_1 , \REG.mem_4_0 , \REG.mem_13_14 , 
        \REG.mem_13_4 , wr_fifo_en_w, rd_fifo_en_w_adj_56, rd_fifo_en_prev_r;
    wire [2:0]wr_addr_r_adj_118;   // src/fifo_quad_word_mod.v(65[31:40])
    wire [2:0]wr_addr_p1_w_adj_120;   // src/fifo_quad_word_mod.v(67[32:44])
    wire [2:0]rd_addr_r_adj_121;   // src/fifo_quad_word_mod.v(69[31:40])
    wire [2:0]rd_addr_p1_w_adj_123;   // src/fifo_quad_word_mod.v(71[32:44])
    
    wire n10871;
    wire [31:0]\mem_LUT.data_raw_r ;   // src/fifo_quad_word_mod.v(449[42:52])
    
    wire empty_o_N_1149, n7473, n6127, n2944, \REG.mem_3_15 , \REG.mem_3_14 , 
        \REG.mem_3_13 , \REG.mem_3_12 , \REG.mem_3_11 , \REG.mem_3_10 , 
        \REG.mem_3_9 , \REG.mem_3_8 , \REG.mem_3_7 , \REG.mem_3_6 , 
        \REG.mem_3_5 , \REG.mem_3_4 , \REG.mem_3_3 , \REG.mem_3_2 , 
        \REG.mem_3_1 , n3022, n4869, n4860, n4859, n6121, n6118, 
        \REG.mem_12_9 , \REG.mem_12_8 , \REG.mem_12_7 , n843, \REG.mem_12_6 , 
        n10430, n6112, n10786, n4459, \REG.mem_12_15 , \REG.mem_12_14 , 
        \REG.mem_12_13 , \REG.mem_12_12 , n10226, \REG.mem_12_11 , \REG.mem_12_10 , 
        \REG.mem_12_4 , \REG.mem_12_5 , n10564, n6106, n1774, n6105, 
        n15, \REG.mem_23_0 , \REG.mem_23_1 , \REG.mem_23_2 , \REG.mem_23_3 , 
        \REG.mem_23_4 , \REG.mem_23_5 , \REG.mem_23_6 , \REG.mem_23_7 , 
        \REG.mem_23_8 , \REG.mem_23_9 , \REG.mem_23_10 , \REG.mem_23_11 , 
        \REG.mem_23_12 , \REG.mem_23_13 , \REG.mem_23_14 , \REG.mem_23_15 , 
        n4192, n14025, \REG.mem_25_0 , \REG.mem_25_1 , \REG.mem_25_2 , 
        \REG.mem_25_3 , \REG.mem_25_4 , \REG.mem_25_5 , \REG.mem_25_6 , 
        \REG.mem_25_7 , \REG.mem_25_8 , \REG.mem_25_9 , \REG.mem_25_10 , 
        \REG.mem_25_11 , \REG.mem_25_12 , \REG.mem_25_13 , \REG.mem_25_14 , 
        \REG.mem_25_15 , n4_adj_58, \REG.mem_31_0 , \REG.mem_31_1 , 
        \REG.mem_31_2 , \REG.mem_31_3 , \REG.mem_31_4 , \REG.mem_31_5 , 
        \REG.mem_31_6 , \REG.mem_31_7 , \REG.mem_31_8 , \REG.mem_31_9 , 
        \REG.mem_31_10 , \REG.mem_31_11 , \REG.mem_31_12 , \REG.mem_31_13 , 
        \REG.mem_31_14 , \REG.mem_31_15 , n10808, \REG.mem_35_0 , \REG.mem_35_1 , 
        \REG.mem_35_2 , \REG.mem_35_3 , \REG.mem_35_4 , \REG.mem_35_5 , 
        \REG.mem_35_6 , \REG.mem_35_7 , \REG.mem_35_8 , \REG.mem_35_9 , 
        \REG.mem_35_10 , \REG.mem_35_11 , \REG.mem_35_12 , \REG.mem_35_13 , 
        \REG.mem_35_14 , \REG.mem_35_15 , n10566, \REG.mem_36_0 , \REG.mem_36_1 , 
        \REG.mem_36_2 , \REG.mem_36_3 , \REG.mem_36_4 , \REG.mem_36_5 , 
        \REG.mem_36_6 , \REG.mem_36_7 , \REG.mem_36_8 , \REG.mem_36_9 , 
        \REG.mem_36_10 , \REG.mem_36_11 , \REG.mem_36_12 , \REG.mem_36_13 , 
        \REG.mem_36_14 , \REG.mem_36_15 , n10913, n10568, \REG.mem_37_0 , 
        \REG.mem_37_1 , \REG.mem_37_2 , \REG.mem_37_3 , \REG.mem_37_4 , 
        \REG.mem_37_5 , \REG.mem_37_6 , \REG.mem_37_7 , \REG.mem_37_8 , 
        \REG.mem_37_9 , \REG.mem_37_10 , \REG.mem_37_11 , \REG.mem_37_12 , 
        \REG.mem_37_13 , \REG.mem_37_14 , \REG.mem_37_15 , n10570, \REG.mem_38_0 , 
        \REG.mem_38_1 , \REG.mem_38_2 , \REG.mem_38_3 , \REG.mem_38_4 , 
        \REG.mem_38_5 , \REG.mem_38_6 , \REG.mem_38_7 , \REG.mem_38_8 , 
        \REG.mem_38_9 , \REG.mem_38_10 , \REG.mem_38_11 , \REG.mem_38_12 , 
        \REG.mem_38_13 , \REG.mem_38_14 , \REG.mem_38_15 , n10572, \REG.mem_39_0 , 
        \REG.mem_39_1 , \REG.mem_39_2 , \REG.mem_39_3 , \REG.mem_39_4 , 
        \REG.mem_39_5 , \REG.mem_39_6 , \REG.mem_39_7 , \REG.mem_39_8 , 
        \REG.mem_39_9 , \REG.mem_39_10 , \REG.mem_39_11 , \REG.mem_39_12 , 
        \REG.mem_39_13 , \REG.mem_39_14 , \REG.mem_39_15 , n32, n10574, 
        \REG.mem_40_0 , \REG.mem_40_1 , \REG.mem_40_2 , \REG.mem_40_3 , 
        \REG.mem_40_4 , \REG.mem_40_5 , \REG.mem_40_6 , \REG.mem_40_7 , 
        \REG.mem_40_8 , \REG.mem_40_9 , \REG.mem_40_10 , \REG.mem_40_11 , 
        \REG.mem_40_12 , \REG.mem_40_13 , \REG.mem_40_14 , \REG.mem_40_15 , 
        \REG.mem_41_0 , \REG.mem_41_1 , \REG.mem_41_2 , \REG.mem_41_3 , 
        \REG.mem_41_4 , \REG.mem_41_5 , \REG.mem_41_6 , \REG.mem_41_7 , 
        \REG.mem_41_8 , \REG.mem_41_9 , \REG.mem_41_10 , \REG.mem_41_11 , 
        \REG.mem_41_12 , \REG.mem_41_13 , \REG.mem_41_14 , \REG.mem_41_15 , 
        n10576, n24, \REG.mem_42_0 , \REG.mem_42_1 , \REG.mem_42_2 , 
        \REG.mem_42_3 , \REG.mem_42_4 , \REG.mem_42_5 , \REG.mem_42_6 , 
        \REG.mem_42_7 , \REG.mem_42_8 , \REG.mem_42_9 , \REG.mem_42_10 , 
        \REG.mem_42_11 , \REG.mem_42_12 , \REG.mem_42_13 , \REG.mem_42_14 , 
        \REG.mem_42_15 , n10578, \REG.mem_43_0 , \REG.mem_43_1 , \REG.mem_43_2 , 
        \REG.mem_43_3 , \REG.mem_43_4 , \REG.mem_43_5 , \REG.mem_43_6 , 
        \REG.mem_43_7 , \REG.mem_43_8 , \REG.mem_43_9 , \REG.mem_43_10 , 
        \REG.mem_43_11 , \REG.mem_43_12 , \REG.mem_43_13 , \REG.mem_43_14 , 
        \REG.mem_43_15 , n6088, \REG.mem_44_0 , \REG.mem_44_1 , \REG.mem_44_2 , 
        \REG.mem_44_3 , \REG.mem_44_4 , \REG.mem_44_5 , \REG.mem_44_6 , 
        \REG.mem_44_7 , \REG.mem_44_8 , \REG.mem_44_9 , \REG.mem_44_10 , 
        \REG.mem_44_11 , \REG.mem_44_12 , \REG.mem_44_13 , \REG.mem_44_14 , 
        \REG.mem_44_15 , \REG.mem_45_0 , \REG.mem_45_1 , \REG.mem_45_2 , 
        \REG.mem_45_3 , \REG.mem_45_4 , \REG.mem_45_5 , \REG.mem_45_6 , 
        \REG.mem_45_7 , \REG.mem_45_8 , \REG.mem_45_9 , \REG.mem_45_10 , 
        \REG.mem_45_11 , \REG.mem_45_12 , \REG.mem_45_13 , \REG.mem_45_14 , 
        \REG.mem_45_15 , \REG.mem_46_0 , \REG.mem_46_1 , \REG.mem_46_2 , 
        \REG.mem_46_3 , \REG.mem_46_4 , \REG.mem_46_5 , \REG.mem_46_6 , 
        \REG.mem_46_7 , \REG.mem_46_8 , \REG.mem_46_9 , \REG.mem_46_10 , 
        \REG.mem_46_11 , \REG.mem_46_12 , \REG.mem_46_13 , \REG.mem_46_14 , 
        \REG.mem_46_15 , n6085, \REG.mem_47_0 , \REG.mem_47_1 , \REG.mem_47_2 , 
        \REG.mem_47_3 , \REG.mem_47_4 , \REG.mem_47_5 , \REG.mem_47_6 , 
        \REG.mem_47_7 , \REG.mem_47_8 , \REG.mem_47_9 , \REG.mem_47_10 , 
        \REG.mem_47_11 , \REG.mem_47_12 , \REG.mem_47_13 , \REG.mem_47_14 , 
        \REG.mem_47_15 , n3495, \REG.mem_48_0 , \REG.mem_48_1 , \REG.mem_48_2 , 
        \REG.mem_48_3 , \REG.mem_48_4 , \REG.mem_48_5 , \REG.mem_48_6 , 
        \REG.mem_48_7 , \REG.mem_48_8 , \REG.mem_48_9 , \REG.mem_48_10 , 
        \REG.mem_48_11 , \REG.mem_48_12 , \REG.mem_48_13 , \REG.mem_48_14 , 
        \REG.mem_48_15 , n6082, n6081, \REG.mem_50_0 , \REG.mem_50_1 , 
        \REG.mem_50_2 , \REG.mem_50_3 , \REG.mem_50_4 , \REG.mem_50_5 , 
        \REG.mem_50_6 , \REG.mem_50_7 , \REG.mem_50_8 , \REG.mem_50_9 , 
        \REG.mem_50_10 , \REG.mem_50_11 , \REG.mem_50_12 , \REG.mem_50_13 , 
        \REG.mem_50_14 , \REG.mem_50_15 , n6079, n10345, n6078, \REG.mem_55_0 , 
        \REG.mem_55_1 , \REG.mem_55_2 , \REG.mem_55_3 , \REG.mem_55_4 , 
        \REG.mem_55_5 , \REG.mem_55_6 , \REG.mem_55_7 , \REG.mem_55_8 , 
        \REG.mem_55_9 , \REG.mem_55_10 , \REG.mem_55_11 , \REG.mem_55_12 , 
        \REG.mem_55_13 , \REG.mem_55_14 , \REG.mem_55_15 , \REG.mem_57_0 , 
        \REG.mem_57_1 , \REG.mem_57_2 , \REG.mem_57_3 , \REG.mem_57_4 , 
        \REG.mem_57_5 , \REG.mem_57_6 , \REG.mem_57_7 , \REG.mem_57_8 , 
        \REG.mem_57_9 , \REG.mem_57_10 , \REG.mem_57_11 , \REG.mem_57_12 , 
        \REG.mem_57_13 , \REG.mem_57_14 , \REG.mem_57_15 , n12063, n10562, 
        n10983, \REG.mem_63_0 , \REG.mem_63_1 , \REG.mem_63_2 , \REG.mem_63_3 , 
        \REG.mem_63_4 , \REG.mem_63_5 , \REG.mem_63_6 , \REG.mem_63_7 , 
        \REG.mem_63_8 , \REG.mem_63_9 , \REG.mem_63_10 , \REG.mem_63_11 , 
        \REG.mem_63_12 , \REG.mem_63_13 , \REG.mem_63_14 , \REG.mem_63_15 , 
        n2, n8_adj_59, n10, n15_adj_60, n17, n18, n19, n20, 
        n21, n22, n23, n24_adj_61, n25, n26, n27, n28, n29, 
        n30, n34, n40, n42, n47, n49, n50, n51, n52, n53, 
        n54, n55, n56, n57, n58, n59, n60, n61, n62, n6077, 
        n6075, n6074, n10580, n10582, n63, n10406, n6060, n6059, 
        n6058, n6057, n6056, n6055, n6054, n6045, n6043, n6024, 
        n6021, n6020, n6019, n6018, n6017, n6016, n6015, n6014, 
        n6013, n6012, n6011, n6010, n6009, n6008, n6007, n6006, 
        n5989, n5970, n5953, n5952, n5951, n5950, n5949, n5948, 
        n5947, n5946, n5945, n5928, n5927, n5926, n5924, n5923, 
        n5921, n5901, n5900, n5899, n5898, n5897, n5896, n5895, 
        n5894, n5893, n5892, n5891, n5890, n5889, n5888, n5887, 
        n5885, n10556, n5868, n5864, n5863, n5862, n5861, n5860, 
        n5859, n5858, n5857, n5856, n5855, n5854, n5853, n5852, 
        n5851, n5850, n5849, n5848, n5847, n5846, n5845, n5844, 
        n5843, n5842, n5841, n5839, n5838, n5837, n5836, n5771, 
        n5770, n5769, n5768, n5767, n5766, n5765, n5764, n5763, 
        n5762, n5761, n5760, n5759, n5758, n5757, n5753, n10514, 
        n5736, n3794, n5735, n5734, n5733, n5732, n5731, n5730, 
        n5729, n5728, n5727, n5726, n5725, n5724, n5723, n5722, 
        n5721, n5720, n5719, n5718, n5717, n5716, n5715, n5714, 
        n5713, n5712, n5711, n5710, n5709, n5708, n5707, n5706, 
        n5705, n5704, n5703, n5702, n5701, n5700, n5699, n5698, 
        n5697, n5696, n5695, n5694, n5693, n5692, n5691, n5690, 
        n5689, n5688, n5687, n5686, n5685, n5684, n5683, n5682, 
        n5681, n5680, n5679, n5678, n5677, n5676, n5675, n5674, 
        n5673, n5671, n5670, n5669, n5668, n5666, n5665, n5664, 
        n5662, n5661, n5660, n5659, n5658, n5657, n5656, n5655, 
        n5654, n5653, n5652, n5651, n5650, n5649, n5648, n5647, 
        n5646, n5645, n5644, n5643, n5642, n5641, n5640, n5639, 
        n5638, n5637, n5636, n5635, n5634, n5633, n5632, n5631, 
        n5630, n5629, n5628, n5627, n5626, n5625, n5624, n5623, 
        n5622, n5621, n5620, n5619, n5618, n5617, n5616, n5615, 
        n5614, n5613, n5612, n5611, n5610, n5609, n5608, n5607, 
        n5606, n5605, n5604, n5603, n5602, n5601, n5600, n5599, 
        n5598, n5597, n5596, n5595, n5594, n5593, n5592, n5591, 
        n5590, n5589, n5588, n5587, n5586, n5585, n5584, n5583, 
        n5582, n5581, n5580, n5579, n5578, n5577, n5576, n5575, 
        n5573, n5572, n5571, n5570, n5569, n5568, n5567, n5566, 
        n5565, n5564, n5563, n5562, n5561, n5560, n5559, n10831, 
        n5558, n5556, n5555, n5554, n5553, n5552, n5551, n5550, 
        n5549, n5548, n5547, n5546, n5545, n5544, n5543, n5542, 
        n5541, n5540, n5539, n5536, n5533, n5532, n5531, n5530, 
        n5529, n5528, n5527, n4248, n5526, n5525, n5524, n5523, 
        n5522, n5521, n5520, n5519, n5518, n5517, n5516, n5515, 
        n5514, n5513, n5512, n5511, n5510, n5507, n5506, n5505, 
        n5504, n5503, n5502, n5501, n5500, n5499, n5498, n5497, 
        n5496, n5495, n10195, n10194, n5494, n5493, n5492, n10193, 
        n10192, n10191, n10190, n10189, n10188, n10187, n130, 
        n129, n128, n127, n126, n125, n124, n123, n122, n121, 
        n120, n5441, n5440, n5439, n5438, n5437, n5436, n5435, 
        n5434, n5433, n5432, n5431, n119, n118, n117, n116, 
        n115, n114, n113, n112, n111, n110, n109, n108, n107, 
        n106, n5430, n5429, n5428, n5427, n5426, n10186, n10185, 
        n10184, n10183, n10182, n10181, n10180, n10179, n10178, 
        n25_adj_62, n24_adj_63, n23_adj_64, n22_adj_65, n21_adj_66, 
        n5345, n5344, n5343, n5342, n5341, n5340, n5339, n5338, 
        n5337, n5336, n5335, n20_adj_67, n19_adj_68, n18_adj_69, 
        n17_adj_70, n16, n15_adj_71, n14, n13, n12, n11, n10_adj_72, 
        n9, n8_adj_73, n7, n6, n5, n5334, n5333, n5332, n5331, 
        n5330, n4_adj_74, n3, n2_adj_75, n10177, n25_adj_76, n5314, 
        n5311, n5306, n5305, n5304, n5303, n5302, n5301, n5300, 
        n5299, n5298, n5297, n5296, n5295, n5294, n5293, n5292, 
        n5290, n4855, n10176, n10175, n10174, n10173, n10172, 
        n10917, n10064, n5224, n5223, n5222, n5221, n5220, n5219, 
        n5218, n5217, n5216, n5215, n5214, n5213, n5212, n5211, 
        n5210, n5209, n4845, n4838, n5192, n5191, n5190, n5189, 
        n5188, n5187, n5186, n5185, n5184, n5183, n5182, n5181, 
        n5180, n5179, n5178, n5177, n5176, n5175, n5174, n5173, 
        n5172, n5171, n5170, n5169, n5168, n5167, n5166, n5165, 
        n5164, n5163, n5162, n5161, n5160, n5159, n5158, n5157, 
        n5156, n5155, n5154, n4824, n5153, n5152, n5151, n5150, 
        n5149, n5148, n5147, n5146, n5145, n5144, n5143, n5142, 
        n5141, n5140, n5139, n5138, n5137, n5136, n5135, n5134, 
        n5133, n5132, n5131, n5130, n5129, n5128, n4836, n4834, 
        n5127, n5126, n5125, n5124, n5123, n5122, n5121, n5120, 
        n5119, n5118, n5117, n5116, n5115, n5114, n5113, n5112, 
        n5111, n5110, n5109, n5108, n5107, n5106, n5105, n5104, 
        n5103, n5102, n5101, n5100, n5099, n5098, n5097, n5096, 
        n5095, n5094, n5093, n5092, n5091, n5090, n5089, n5088, 
        n5087, n5086, n5085, n5084, n5083, n5082, n5081, n5080, 
        n5079, n5078, n5077, n5076, n5075, n5074, n5073, n5072, 
        n5071, n5070, n5069, n5068, n5067, n5066, n5065, n5064, 
        n5063, n5062, n5061, n5060, n5059, n5057, n5056, n5055, 
        n5054, n5053, n5052, n5051, n5050, n5049, n5048, n5047, 
        n5046, n5045, n5044, n5043, n5042, n5041, n5040, n5039, 
        n5038, n5037, n5036, n5035, n5034, n5033, n5032, n5031, 
        n5030, n5029, n5028, n5027, n5026, n5025, n5024, n5023, 
        n5022, n5021, n5020, n5019, n5018, n5017, n5016, n5015, 
        n10897, n10877, n10873, n5014, n5013, n5012, n5011, n5010, 
        n5009, n5008, n5007, n5006, n5005, n10805, n5004, n5003, 
        n5002, n5001, n5000, n4999, n4998, n4997, n4996, n4995, 
        n4994, n4993, n4992, n4991, n4990, n4989, n4988, n4987, 
        n4986, n4985, n4984, n4983, n4982, n4981, n4980, n4979, 
        n4335, n4978, n4977, n4976, n4319, n4975, n4974, n4973, 
        n4972, n4312, n4_adj_77, n4971, n4970, n4_adj_78, n4969, 
        n4968, n4967, n4966, n4965, n4964, n4963, n4962, n4961, 
        n10295, n1, n10588, n13865, n10293, n10291;
    
    VCC i2 (.Y(VCC_net));
    timing_controller timing_controller_inst (.state({state}), .SLM_CLK_c(SLM_CLK_c), 
            .n1879(n1879), .GND_net(GND_net), .n10514(n10514), .VCC_net(VCC_net), 
            .n10808(n10808), .reset_per_frame(reset_per_frame), .n1774(n1774), 
            .n7386(n7386), .INVERT_c_3(INVERT_c_3), .buffer_switch_done(buffer_switch_done), 
            .n4245(n4245), .n7568(n7568), .n7590(n7590), .n4192(n4192), 
            .n63(n63), .n10831(n10831), .UPDATE_c_2(UPDATE_c_2)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(452[19] 464[2])
    SB_LUT4 i4623_3_lut (.I0(\REG.mem_63_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n2), .I3(GND_net), .O(n6006));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4127_3_lut (.I0(tx_data_byte[6]), .I1(pc_data_rx[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5510));   // src/top.v(1074[8] 1141[4])
    defparam i4127_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF uart_rx_complete_prev_83 (.Q(uart_rx_complete_prev), .C(SLM_CLK_c), 
           .D(debug_led3));   // src/top.v(1065[8] 1071[4])
    bluejay_data bluejay_data_inst (.dc32_fifo_almost_full(dc32_fifo_almost_full), 
            .n771(n771), .dc32_fifo_almost_empty(dc32_fifo_almost_empty), 
            .bluejay_data_out_31__N_736(bluejay_data_out_31__N_736), .buffer_switch_done_latched(buffer_switch_done_latched), 
            .GND_net(GND_net), .DEBUG_9_c(DEBUG_9_c), .SLM_CLK_c(SLM_CLK_c), 
            .DATA19_c(DATA19_c), .buffer_switch_done(buffer_switch_done), 
            .n4937(n4937), .DATA18_c(DATA18_c), .n4936(n4936), .DATA17_c(DATA17_c), 
            .n6112(n6112), .DEBUG_6_c(DEBUG_6_c), .DATA15_c(DATA15_c), 
            .DATA14_c(DATA14_c), .DATA13_c(DATA13_c), .DATA12_c(DATA12_c), 
            .n843(n843), .VCC_net(VCC_net), .DATA11_c(DATA11_c), .DATA10_c(DATA10_c), 
            .SYNC_c(SYNC_c), .bluejay_data_out_31__N_737(bluejay_data_out_31__N_737), 
            .n10277(n10277), .DATA9_c(DATA9_c), .DATA8_c(DATA8_c), .DATA7_c(DATA7_c), 
            .DATA6_c(DATA6_c), .\rd_sig_diff0_w[1] (rd_sig_diff0_w[1]), 
            .get_next_word(get_next_word), .\rd_sig_diff0_w[0] (rd_sig_diff0_w[0]), 
            .\rd_sig_diff0_w[2] (rd_sig_diff0_w[2]), .n10873(n10873), .n10877(n10877), 
            .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .DATA5_c(DATA5_c), .DATA20_c(DATA20_c), .\fifo_data_out[4] (fifo_data_out[4]), 
            .\fifo_data_out[5] (fifo_data_out[5]), .\fifo_data_out[6] (fifo_data_out[6]), 
            .\fifo_data_out[7] (fifo_data_out[7]), .\fifo_data_out[11] (fifo_data_out[11]), 
            .\fifo_data_out[10] (fifo_data_out[10]), .\fifo_data_out[3] (fifo_data_out[3]), 
            .\fifo_data_out[15] (fifo_data_out[15]), .\fifo_data_out[14] (fifo_data_out[14]), 
            .\fifo_data_out[13] (fifo_data_out[13]), .\fifo_data_out[12] (fifo_data_out[12]), 
            .\fifo_data_out[9] (fifo_data_out[9]), .\fifo_data_out[8] (fifo_data_out[8])) /* synthesis syn_module_defined=1 */ ;   // src/top.v(626[14] 639[2])
    SB_LUT4 i4128_3_lut (.I0(\REG.mem_36_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n29), .I3(GND_net), .O(n5511));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4128_3_lut.LUT_INIT = 16'hcaca;
    SB_GB clk_gb (.GLOBAL_BUFFER_OUTPUT(SLM_CLK_c), .USER_SIGNAL_TO_GLOBAL_BUFFER(pll_clk_unbuf)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=222, LSE_RLINE=228 */ ;   // src/clock.v(82[7:96])
    SB_LUT4 i4129_3_lut (.I0(\REG.mem_36_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n29), .I3(GND_net), .O(n5512));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4130_3_lut (.I0(\REG.mem_36_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n29), .I3(GND_net), .O(n5513));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4131_3_lut (.I0(\REG.mem_36_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n29), .I3(GND_net), .O(n5514));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4131_3_lut.LUT_INIT = 16'hcaca;
    SB_IO RST_pad (.PACKAGE_PIN(RST), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RST_pad.PIN_TYPE = 6'b011001;
    defparam RST_pad.PULLUP = 1'b0;
    defparam RST_pad.NEG_TRIGGER = 1'b0;
    defparam RST_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i3515_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4898));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i3515_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4624_3_lut (.I0(\REG.mem_63_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n2), .I3(GND_net), .O(n6007));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4625_3_lut (.I0(\REG.mem_63_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n2), .I3(GND_net), .O(n6008));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4132_3_lut (.I0(\REG.mem_36_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n29), .I3(GND_net), .O(n5515));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4133_3_lut (.I0(\REG.mem_36_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n29), .I3(GND_net), .O(n5516));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4134_3_lut (.I0(\REG.mem_36_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n29), .I3(GND_net), .O(n5517));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4135_3_lut (.I0(\REG.mem_36_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n29), .I3(GND_net), .O(n5518));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4626_3_lut (.I0(\REG.mem_63_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n2), .I3(GND_net), .O(n6009));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4627_3_lut (.I0(\REG.mem_63_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n2), .I3(GND_net), .O(n6010));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4136_3_lut (.I0(\REG.mem_36_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n29), .I3(GND_net), .O(n5519));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4137_3_lut (.I0(\REG.mem_36_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n29), .I3(GND_net), .O(n5520));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4198_3_lut (.I0(\REG.mem_39_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n26), .I3(GND_net), .O(n5581));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4138_3_lut (.I0(\REG.mem_36_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n29), .I3(GND_net), .O(n5521));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4139_3_lut (.I0(\REG.mem_36_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n29), .I3(GND_net), .O(n5522));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4199_3_lut (.I0(\REG.mem_39_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n26), .I3(GND_net), .O(n5582));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4140_3_lut (.I0(\REG.mem_36_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n29), .I3(GND_net), .O(n5523));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4141_3_lut (.I0(\REG.mem_36_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n29), .I3(GND_net), .O(n5524));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4141_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_all_r_77 (.Q(reset_all_w), .C(SLM_CLK_c), .D(reset_all_w_N_61));   // src/top.v(246[8] 264[4])
    SB_LUT4 i4200_3_lut (.I0(\REG.mem_39_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n26), .I3(GND_net), .O(n5583));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4142_3_lut (.I0(\REG.mem_36_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n29), .I3(GND_net), .O(n5525));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4143_3_lut (.I0(\REG.mem_36_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n29), .I3(GND_net), .O(n5526));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4144_3_lut (.I0(tx_addr_byte[7]), .I1(tx_data_byte[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5527));   // src/top.v(1074[8] 1141[4])
    defparam i4144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4201_3_lut (.I0(\REG.mem_39_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n26), .I3(GND_net), .O(n5584));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4145_3_lut (.I0(tx_addr_byte[6]), .I1(tx_data_byte[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5528));   // src/top.v(1074[8] 1141[4])
    defparam i4145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4628_3_lut (.I0(\REG.mem_63_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n2), .I3(GND_net), .O(n6011));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4202_3_lut (.I0(\REG.mem_39_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n26), .I3(GND_net), .O(n5585));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4146_3_lut (.I0(tx_addr_byte[5]), .I1(tx_data_byte[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5529));   // src/top.v(1074[8] 1141[4])
    defparam i4146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4203_3_lut (.I0(\REG.mem_39_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n26), .I3(GND_net), .O(n5586));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4147_3_lut (.I0(tx_addr_byte[4]), .I1(tx_data_byte[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5530));   // src/top.v(1074[8] 1141[4])
    defparam i4147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4148_3_lut (.I0(tx_addr_byte[3]), .I1(tx_data_byte[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5531));   // src/top.v(1074[8] 1141[4])
    defparam i4148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4149_3_lut (.I0(tx_addr_byte[2]), .I1(tx_data_byte[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5532));   // src/top.v(1074[8] 1141[4])
    defparam i4149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4204_3_lut (.I0(\REG.mem_39_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n26), .I3(GND_net), .O(n5587));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4205_3_lut (.I0(\REG.mem_39_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n26), .I3(GND_net), .O(n5588));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4629_3_lut (.I0(\REG.mem_63_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n2), .I3(GND_net), .O(n6012));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4630_3_lut (.I0(\REG.mem_63_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n2), .I3(GND_net), .O(n6013));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4631_3_lut (.I0(\REG.mem_63_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n2), .I3(GND_net), .O(n6014));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4150_3_lut (.I0(tx_addr_byte[1]), .I1(tx_data_byte[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5533));   // src/top.v(1074[8] 1141[4])
    defparam i4150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4157_3_lut (.I0(\REG.mem_37_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n28), .I3(GND_net), .O(n5540));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4632_3_lut (.I0(\REG.mem_63_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n2), .I3(GND_net), .O(n6015));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4158_3_lut (.I0(\REG.mem_37_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n28), .I3(GND_net), .O(n5541));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4159_3_lut (.I0(\REG.mem_37_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n28), .I3(GND_net), .O(n5542));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4160_3_lut (.I0(\REG.mem_37_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n28), .I3(GND_net), .O(n5543));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4161_3_lut (.I0(\REG.mem_37_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n28), .I3(GND_net), .O(n5544));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4162_3_lut (.I0(\REG.mem_37_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n28), .I3(GND_net), .O(n5545));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4163_3_lut (.I0(\REG.mem_37_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n28), .I3(GND_net), .O(n5546));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4164_3_lut (.I0(\REG.mem_37_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n28), .I3(GND_net), .O(n5547));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4165_3_lut (.I0(\REG.mem_37_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n28), .I3(GND_net), .O(n5548));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4633_3_lut (.I0(\REG.mem_63_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n2), .I3(GND_net), .O(n6016));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4206_3_lut (.I0(\REG.mem_39_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n26), .I3(GND_net), .O(n5589));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [13]), .I3(fifo_data_out[13]), .O(n10580));
    defparam i12_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4634_3_lut (.I0(\REG.mem_63_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n2), .I3(GND_net), .O(n6017));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4166_3_lut (.I0(\REG.mem_37_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n28), .I3(GND_net), .O(n5549));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4167_3_lut (.I0(\REG.mem_37_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n28), .I3(GND_net), .O(n5550));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4168_3_lut (.I0(\REG.mem_37_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n28), .I3(GND_net), .O(n5551));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4278_3_lut (.I0(\REG.mem_44_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n21), .I3(GND_net), .O(n5661));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4207_3_lut (.I0(\REG.mem_40_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n25), .I3(GND_net), .O(n5590));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4169_3_lut (.I0(\REG.mem_37_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n28), .I3(GND_net), .O(n5552));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4279_3_lut (.I0(\REG.mem_44_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n21), .I3(GND_net), .O(n5662));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4170_3_lut (.I0(\REG.mem_37_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n28), .I3(GND_net), .O(n5553));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4171_3_lut (.I0(\REG.mem_37_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n28), .I3(GND_net), .O(n5554));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4208_3_lut (.I0(\REG.mem_40_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n25), .I3(GND_net), .O(n5591));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4172_3_lut (.I0(\REG.mem_37_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n28), .I3(GND_net), .O(n5555));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4173_3_lut (.I0(\REG.mem_38_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n27), .I3(GND_net), .O(n5556));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4175_3_lut (.I0(\REG.mem_38_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n27), .I3(GND_net), .O(n5558));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4176_3_lut (.I0(\REG.mem_38_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n27), .I3(GND_net), .O(n5559));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4177_3_lut (.I0(\REG.mem_38_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n27), .I3(GND_net), .O(n5560));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_74 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [14]), .I3(fifo_data_out[14]), .O(n10582));
    defparam i12_4_lut_4_lut_adj_74.LUT_INIT = 16'h3120;
    SB_LUT4 i4178_3_lut (.I0(\REG.mem_38_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n27), .I3(GND_net), .O(n5561));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4179_3_lut (.I0(\REG.mem_38_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n27), .I3(GND_net), .O(n5562));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4180_3_lut (.I0(\REG.mem_38_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n27), .I3(GND_net), .O(n5563));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4181_3_lut (.I0(\REG.mem_38_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n27), .I3(GND_net), .O(n5564));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4182_3_lut (.I0(\REG.mem_38_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n27), .I3(GND_net), .O(n5565));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4183_3_lut (.I0(\REG.mem_38_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n27), .I3(GND_net), .O(n5566));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4184_3_lut (.I0(\REG.mem_38_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n27), .I3(GND_net), .O(n5567));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4209_3_lut (.I0(\REG.mem_40_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n25), .I3(GND_net), .O(n5592));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4185_3_lut (.I0(\REG.mem_38_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n27), .I3(GND_net), .O(n5568));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4186_3_lut (.I0(\REG.mem_38_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n27), .I3(GND_net), .O(n5569));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4281_3_lut (.I0(\REG.mem_44_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n21), .I3(GND_net), .O(n5664));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4282_3_lut (.I0(\REG.mem_44_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n21), .I3(GND_net), .O(n5665));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4210_3_lut (.I0(\REG.mem_40_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n25), .I3(GND_net), .O(n5593));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4187_3_lut (.I0(\REG.mem_38_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n27), .I3(GND_net), .O(n5570));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4211_3_lut (.I0(\REG.mem_40_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n25), .I3(GND_net), .O(n5594));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4212_3_lut (.I0(\REG.mem_40_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n25), .I3(GND_net), .O(n5595));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4188_3_lut (.I0(\REG.mem_38_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n27), .I3(GND_net), .O(n5571));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_75 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [12]), .I3(fifo_data_out[12]), .O(n10578));
    defparam i12_4_lut_4_lut_adj_75.LUT_INIT = 16'h3120;
    SB_LUT4 i4283_3_lut (.I0(\REG.mem_44_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n21), .I3(GND_net), .O(n5666));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4635_3_lut (.I0(\REG.mem_63_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n2), .I3(GND_net), .O(n6018));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4189_3_lut (.I0(\REG.mem_38_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n27), .I3(GND_net), .O(n5572));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4285_3_lut (.I0(\REG.mem_44_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n21), .I3(GND_net), .O(n5668));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4190_3_lut (.I0(\REG.mem_39_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n26), .I3(GND_net), .O(n5573));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4286_3_lut (.I0(\REG.mem_44_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n21), .I3(GND_net), .O(n5669));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4702_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [0]), .I3(fifo_data_out[0]), .O(n6085));
    defparam i4702_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4287_3_lut (.I0(\REG.mem_44_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n21), .I3(GND_net), .O(n5670));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4636_3_lut (.I0(\REG.mem_63_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n2), .I3(GND_net), .O(n6019));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4213_3_lut (.I0(\REG.mem_40_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n25), .I3(GND_net), .O(n5596));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4192_3_lut (.I0(\REG.mem_39_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n26), .I3(GND_net), .O(n5575));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4193_3_lut (.I0(\REG.mem_39_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n26), .I3(GND_net), .O(n5576));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_76 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [11]), .I3(fifo_data_out[11]), .O(n10576));
    defparam i12_4_lut_4_lut_adj_76.LUT_INIT = 16'h3120;
    SB_LUT4 i4194_3_lut (.I0(\REG.mem_39_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n26), .I3(GND_net), .O(n5577));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3516_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4899));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i3516_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4195_3_lut (.I0(\REG.mem_39_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n26), .I3(GND_net), .O(n5578));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4196_3_lut (.I0(\REG.mem_39_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n26), .I3(GND_net), .O(n5579));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4197_3_lut (.I0(\REG.mem_39_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n26), .I3(GND_net), .O(n5580));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3514_3_lut (.I0(rx_buf_byte[0]), .I1(rx_shift_reg[0]), .I2(n3495), 
            .I3(GND_net), .O(n4897));   // src/spi.v(76[8] 221[4])
    defparam i3514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4288_3_lut (.I0(\REG.mem_44_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n21), .I3(GND_net), .O(n5671));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_77 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [10]), .I3(fifo_data_out[10]), .O(n10574));
    defparam i12_4_lut_4_lut_adj_77.LUT_INIT = 16'h3120;
    SB_LUT4 i4738_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [2]), .I3(fifo_data_out[2]), .O(n6121));
    defparam i4738_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4637_3_lut (.I0(\REG.mem_63_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n2), .I3(GND_net), .O(n6020));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4290_3_lut (.I0(\REG.mem_45_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n20), .I3(GND_net), .O(n5673));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4291_3_lut (.I0(\REG.mem_45_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n20), .I3(GND_net), .O(n5674));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4292_3_lut (.I0(\REG.mem_45_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n20), .I3(GND_net), .O(n5675));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3539_4_lut (.I0(RESET_c), .I1(rd_addr_r_adj_121[2]), .I2(rd_addr_p1_w_adj_123[2]), 
            .I3(empty_o_N_1149), .O(n4922));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i3539_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i4109_3_lut (.I0(\REG.mem_35_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n30), .I3(GND_net), .O(n5492));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4293_3_lut (.I0(\REG.mem_45_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n20), .I3(GND_net), .O(n5676));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3520_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4903));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i3520_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4110_3_lut (.I0(\REG.mem_35_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n30), .I3(GND_net), .O(n5493));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4294_3_lut (.I0(\REG.mem_45_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n20), .I3(GND_net), .O(n5677));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3521_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4904));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i3521_2_lut.LUT_INIT = 16'h4444;
    SB_DFF tx_data_byte_r_i0_i7 (.Q(tx_data_byte[7]), .C(SLM_CLK_c), .D(n4942));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 i3524_2_lut (.I0(n2352), .I1(DEBUG_8_c_0_c), .I2(GND_net), 
            .I3(GND_net), .O(n4907));   // src/usb3_if.v(88[8] 191[4])
    defparam i3524_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3526_2_lut (.I0(uart_rx_complete_prev), .I1(debug_led3), .I2(GND_net), 
            .I3(GND_net), .O(n4909));   // src/top.v(1065[8] 1071[4])
    defparam i3526_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3527_2_lut (.I0(reset_per_frame_latched), .I1(n571), .I2(GND_net), 
            .I3(GND_net), .O(n4910));   // src/usb3_if.v(98[9] 189[16])
    defparam i3527_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4295_3_lut (.I0(\REG.mem_45_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n20), .I3(GND_net), .O(n5678));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4214_3_lut (.I0(\REG.mem_40_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n25), .I3(GND_net), .O(n5597));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4638_3_lut (.I0(\REG.mem_63_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n2), .I3(GND_net), .O(n6021));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4111_3_lut (.I0(\REG.mem_35_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n30), .I3(GND_net), .O(n5494));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4215_3_lut (.I0(\REG.mem_40_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n25), .I3(GND_net), .O(n5598));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4215_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF fifo_write_cmd_79 (.Q(fifo_write_cmd), .C(SLM_CLK_c), .D(n4939));   // src/top.v(889[8] 898[4])
    SB_LUT4 i4216_3_lut (.I0(\REG.mem_40_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n25), .I3(GND_net), .O(n5599));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_78 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [15]), .I3(fifo_data_out[15]), .O(n10588));
    defparam i12_4_lut_4_lut_adj_78.LUT_INIT = 16'h3120;
    SB_LUT4 i4112_3_lut (.I0(\REG.mem_35_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n30), .I3(GND_net), .O(n5495));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4217_3_lut (.I0(\REG.mem_40_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n25), .I3(GND_net), .O(n5600));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4113_3_lut (.I0(\REG.mem_35_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n30), .I3(GND_net), .O(n5496));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4296_3_lut (.I0(\REG.mem_45_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n20), .I3(GND_net), .O(n5679));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4297_3_lut (.I0(\REG.mem_45_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n20), .I3(GND_net), .O(n5680));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4114_3_lut (.I0(\REG.mem_35_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n30), .I3(GND_net), .O(n5497));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4218_3_lut (.I0(\REG.mem_40_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n25), .I3(GND_net), .O(n5601));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4115_3_lut (.I0(\REG.mem_35_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n30), .I3(GND_net), .O(n5498));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4298_3_lut (.I0(\REG.mem_45_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n20), .I3(GND_net), .O(n5681));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4219_3_lut (.I0(\REG.mem_40_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n25), .I3(GND_net), .O(n5602));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4219_3_lut.LUT_INIT = 16'hcaca;
    SB_IO CTS_pad (.PACKAGE_PIN(CTS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CTS_pad.PIN_TYPE = 6'b011001;
    defparam CTS_pad.PULLUP = 1'b0;
    defparam CTS_pad.NEG_TRIGGER = 1'b0;
    defparam CTS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY led_counter_1186_1260_add_4_6 (.CI(n10175), .I0(GND_net), .I1(n21_adj_66), 
            .CO(n10176));
    SB_LUT4 i4299_3_lut (.I0(\REG.mem_45_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n20), .I3(GND_net), .O(n5682));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4299_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DTR_pad (.PACKAGE_PIN(DTR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DTR_pad.PIN_TYPE = 6'b011001;
    defparam DTR_pad.PULLUP = 1'b0;
    defparam DTR_pad.NEG_TRIGGER = 1'b0;
    defparam DTR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4116_3_lut (.I0(\REG.mem_35_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n30), .I3(GND_net), .O(n5499));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4116_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DSR_pad (.PACKAGE_PIN(DSR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DSR_pad.PIN_TYPE = 6'b011001;
    defparam DSR_pad.PULLUP = 1'b0;
    defparam DSR_pad.NEG_TRIGGER = 1'b0;
    defparam DSR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4117_3_lut (.I0(\REG.mem_35_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n30), .I3(GND_net), .O(n5500));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4117_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DCD_pad (.PACKAGE_PIN(DCD), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DCD_pad.PIN_TYPE = 6'b011001;
    defparam DCD_pad.PULLUP = 1'b0;
    defparam DCD_pad.NEG_TRIGGER = 1'b0;
    defparam DCD_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4118_3_lut (.I0(\REG.mem_35_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n30), .I3(GND_net), .O(n5501));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4118_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DEBUG_8_c_0_pad (.PACKAGE_PIN(FIFO_D0), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(DEBUG_8_c_0_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_8_c_0_pad.PIN_TYPE = 6'b000001;
    defparam DEBUG_8_c_0_pad.PULLUP = 1'b0;
    defparam DEBUG_8_c_0_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_8_c_0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4220_3_lut (.I0(\REG.mem_40_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n25), .I3(GND_net), .O(n5603));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4221_3_lut (.I0(\REG.mem_40_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n25), .I3(GND_net), .O(n5604));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_79 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [4]), .I3(fifo_data_out[4]), .O(n10562));
    defparam i12_4_lut_4_lut_adj_79.LUT_INIT = 16'h3120;
    SB_LUT4 i4300_3_lut (.I0(\REG.mem_45_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n20), .I3(GND_net), .O(n5683));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4301_3_lut (.I0(\REG.mem_45_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n20), .I3(GND_net), .O(n5684));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4119_3_lut (.I0(\REG.mem_35_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n30), .I3(GND_net), .O(n5502));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4302_3_lut (.I0(\REG.mem_45_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n20), .I3(GND_net), .O(n5685));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4641_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[5]), .I2(GND_net), 
            .I3(GND_net), .O(n6024));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4641_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4303_3_lut (.I0(\REG.mem_45_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n20), .I3(GND_net), .O(n5686));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4222_3_lut (.I0(\REG.mem_40_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n25), .I3(GND_net), .O(n5605));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4223_3_lut (.I0(\REG.mem_41_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5606));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_80 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [8]), .I3(fifo_data_out[8]), .O(n10570));
    defparam i12_4_lut_4_lut_adj_80.LUT_INIT = 16'h3120;
    SB_LUT4 i4304_3_lut (.I0(\REG.mem_45_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n20), .I3(GND_net), .O(n5687));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4224_3_lut (.I0(\REG.mem_41_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5607));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4225_3_lut (.I0(\REG.mem_41_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5608));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_81 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [6]), .I3(fifo_data_out[6]), .O(n10566));
    defparam i12_4_lut_4_lut_adj_81.LUT_INIT = 16'h3120;
    SB_LUT4 i4120_3_lut (.I0(\REG.mem_35_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n30), .I3(GND_net), .O(n5503));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4305_3_lut (.I0(\REG.mem_45_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n20), .I3(GND_net), .O(n5688));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4735_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [1]), .I3(fifo_data_out[1]), .O(n6118));
    defparam i4735_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4306_3_lut (.I0(\REG.mem_46_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n19), .I3(GND_net), .O(n5689));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4226_3_lut (.I0(\REG.mem_41_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5609));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4307_3_lut (.I0(\REG.mem_46_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n19), .I3(GND_net), .O(n5690));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_82 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [7]), .I3(fifo_data_out[7]), .O(n10568));
    defparam i12_4_lut_4_lut_adj_82.LUT_INIT = 16'h3120;
    SB_LUT4 i4227_3_lut (.I0(\REG.mem_41_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5610));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4228_3_lut (.I0(\REG.mem_41_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5611));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4308_3_lut (.I0(\REG.mem_46_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n19), .I3(GND_net), .O(n5691));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4309_3_lut (.I0(\REG.mem_46_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n19), .I3(GND_net), .O(n5692));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4121_3_lut (.I0(\REG.mem_35_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n30), .I3(GND_net), .O(n5504));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4122_3_lut (.I0(\REG.mem_35_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n30), .I3(GND_net), .O(n5505));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4310_3_lut (.I0(\REG.mem_46_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n19), .I3(GND_net), .O(n5693));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3528_2_lut (.I0(reset_per_frame_latched), .I1(n575), .I2(GND_net), 
            .I3(GND_net), .O(n4911));   // src/usb3_if.v(98[9] 189[16])
    defparam i3528_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4123_3_lut (.I0(\REG.mem_35_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n30), .I3(GND_net), .O(n5506));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4229_3_lut (.I0(\REG.mem_41_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5612));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4311_3_lut (.I0(\REG.mem_46_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n19), .I3(GND_net), .O(n5694));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4312_3_lut (.I0(\REG.mem_46_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n19), .I3(GND_net), .O(n5695));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4313_3_lut (.I0(\REG.mem_46_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n19), .I3(GND_net), .O(n5696));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4314_3_lut (.I0(\REG.mem_46_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n19), .I3(GND_net), .O(n5697));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4314_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i0 (.Q(n25_adj_62), .C(SLM_CLK_c), .D(n130));   // src/top.v(203[20:35])
    SB_LUT4 i4315_3_lut (.I0(\REG.mem_46_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n19), .I3(GND_net), .O(n5698));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_83 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [3]), .I3(fifo_data_out[3]), .O(n10556));
    defparam i12_4_lut_4_lut_adj_83.LUT_INIT = 16'h3120;
    SB_LUT4 i4316_3_lut (.I0(\REG.mem_46_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n19), .I3(GND_net), .O(n5699));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_84 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [5]), .I3(fifo_data_out[5]), .O(n10564));
    defparam i12_4_lut_4_lut_adj_84.LUT_INIT = 16'h3120;
    SB_LUT4 i4124_3_lut (.I0(\REG.mem_35_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n30), .I3(GND_net), .O(n5507));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4317_3_lut (.I0(\REG.mem_46_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n19), .I3(GND_net), .O(n5700));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4318_3_lut (.I0(\REG.mem_46_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n19), .I3(GND_net), .O(n5701));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4318_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_clk_counter_i3_1187__i3 (.Q(reset_clk_counter[3]), .C(SLM_CLK_c), 
           .D(n10293));   // src/top.v(259[27:51])
    SB_LUT4 i12_4_lut_4_lut_adj_85 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [9]), .I3(fifo_data_out[9]), .O(n10572));
    defparam i12_4_lut_4_lut_adj_85.LUT_INIT = 16'h3120;
    SB_LUT4 i4230_3_lut (.I0(\REG.mem_41_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5613));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4319_3_lut (.I0(\REG.mem_46_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n19), .I3(GND_net), .O(n5702));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4231_3_lut (.I0(\REG.mem_41_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5614));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4232_3_lut (.I0(\REG.mem_41_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5615));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3540_3_lut (.I0(tx_addr_byte[0]), .I1(tx_data_byte[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4923));   // src/top.v(1074[8] 1141[4])
    defparam i3540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4233_3_lut (.I0(\REG.mem_41_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5616));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4234_3_lut (.I0(\REG.mem_41_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5617));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4320_3_lut (.I0(\REG.mem_46_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n19), .I3(GND_net), .O(n5703));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4235_3_lut (.I0(\REG.mem_41_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5618));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4321_3_lut (.I0(\REG.mem_46_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n19), .I3(GND_net), .O(n5704));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4321_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_clk_counter_i3_1187__i2 (.Q(reset_clk_counter[2]), .C(SLM_CLK_c), 
           .D(n10295));   // src/top.v(259[27:51])
    SB_DFF reset_clk_counter_i3_1187__i1 (.Q(reset_clk_counter[1]), .C(SLM_CLK_c), 
           .D(n10291));   // src/top.v(259[27:51])
    SB_DFF led_counter_1186_1260__i24 (.Q(DEBUG_0_c_24), .C(SLM_CLK_c), 
           .D(n106));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i23 (.Q(n2_adj_75), .C(SLM_CLK_c), .D(n107));   // src/top.v(203[20:35])
    SB_LUT4 i4236_3_lut (.I0(\REG.mem_41_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5619));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4236_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i22 (.Q(n3), .C(SLM_CLK_c), .D(n108));   // src/top.v(203[20:35])
    SB_LUT4 i4237_3_lut (.I0(\REG.mem_41_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5620));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4237_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i21 (.Q(n4_adj_74), .C(SLM_CLK_c), .D(n109));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i20 (.Q(n5), .C(SLM_CLK_c), .D(n110));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i19 (.Q(n6), .C(SLM_CLK_c), .D(n111));   // src/top.v(203[20:35])
    SB_LUT4 i4322_3_lut (.I0(\REG.mem_47_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n18), .I3(GND_net), .O(n5705));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4323_3_lut (.I0(\REG.mem_47_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n18), .I3(GND_net), .O(n5706));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4324_3_lut (.I0(\REG.mem_47_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n18), .I3(GND_net), .O(n5707));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4238_3_lut (.I0(\REG.mem_41_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5621));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4325_3_lut (.I0(\REG.mem_47_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n18), .I3(GND_net), .O(n5708));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4239_3_lut (.I0(\REG.mem_42_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n23), .I3(GND_net), .O(n5622));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4326_3_lut (.I0(\REG.mem_47_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n18), .I3(GND_net), .O(n5709));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4326_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i18 (.Q(n7), .C(SLM_CLK_c), .D(n112));   // src/top.v(203[20:35])
    SB_LUT4 i4240_3_lut (.I0(\REG.mem_42_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n23), .I3(GND_net), .O(n5623));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4240_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i17 (.Q(n8_adj_73), .C(SLM_CLK_c), .D(n113));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i16 (.Q(n9), .C(SLM_CLK_c), .D(n114));   // src/top.v(203[20:35])
    SB_LUT4 i4241_3_lut (.I0(\REG.mem_42_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n23), .I3(GND_net), .O(n5624));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4241_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i15 (.Q(n10_adj_72), .C(SLM_CLK_c), .D(n115));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i14 (.Q(n11), .C(SLM_CLK_c), .D(n116));   // src/top.v(203[20:35])
    SB_LUT4 i4327_3_lut (.I0(\REG.mem_47_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n18), .I3(GND_net), .O(n5710));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4327_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i13 (.Q(n12), .C(SLM_CLK_c), .D(n117));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i12 (.Q(n13), .C(SLM_CLK_c), .D(n118));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i11 (.Q(n14), .C(SLM_CLK_c), .D(n119));   // src/top.v(203[20:35])
    SB_LUT4 i4242_3_lut (.I0(\REG.mem_42_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n23), .I3(GND_net), .O(n5625));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4242_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i10 (.Q(n15_adj_71), .C(SLM_CLK_c), .D(n120));   // src/top.v(203[20:35])
    SB_LUT4 i4243_3_lut (.I0(\REG.mem_42_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n23), .I3(GND_net), .O(n5626));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4243_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i9 (.Q(n16), .C(SLM_CLK_c), .D(n121));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i8 (.Q(n17_adj_70), .C(SLM_CLK_c), .D(n122));   // src/top.v(203[20:35])
    SB_LUT4 i4328_3_lut (.I0(\REG.mem_47_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n18), .I3(GND_net), .O(n5711));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4328_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i7 (.Q(n18_adj_69), .C(SLM_CLK_c), .D(n123));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i6 (.Q(n19_adj_68), .C(SLM_CLK_c), .D(n124));   // src/top.v(203[20:35])
    SB_LUT4 i4329_3_lut (.I0(\REG.mem_47_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n18), .I3(GND_net), .O(n5712));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4329_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i5 (.Q(n20_adj_67), .C(SLM_CLK_c), .D(n125));   // src/top.v(203[20:35])
    SB_LUT4 i4244_3_lut (.I0(\REG.mem_42_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n23), .I3(GND_net), .O(n5627));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4244_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i4 (.Q(n21_adj_66), .C(SLM_CLK_c), .D(n126));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i3 (.Q(n22_adj_65), .C(SLM_CLK_c), .D(n127));   // src/top.v(203[20:35])
    SB_LUT4 i4330_3_lut (.I0(\REG.mem_47_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n18), .I3(GND_net), .O(n5713));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4331_3_lut (.I0(\REG.mem_47_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n18), .I3(GND_net), .O(n5714));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_765[2]), 
            .I3(r_SM_Main[0]), .O(n4335));   // src/uart_rx.v(49[10] 144[8])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i4245_3_lut (.I0(\REG.mem_42_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n23), .I3(GND_net), .O(n5628));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4332_3_lut (.I0(\REG.mem_47_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n18), .I3(GND_net), .O(n5715));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4333_3_lut (.I0(\REG.mem_47_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n18), .I3(GND_net), .O(n5716));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4660_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[3]), .I2(GND_net), 
            .I3(GND_net), .O(n6043));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4660_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4334_3_lut (.I0(\REG.mem_47_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n18), .I3(GND_net), .O(n5717));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4334_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i2 (.Q(n23_adj_64), .C(SLM_CLK_c), .D(n128));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i1 (.Q(n24_adj_63), .C(SLM_CLK_c), .D(n129));   // src/top.v(203[20:35])
    SB_LUT4 i1_4_lut (.I0(rd_addr_r_adj_121[1]), .I1(rd_addr_r_adj_121[0]), 
            .I2(wr_addr_r_adj_118[1]), .I3(wr_addr_r_adj_118[0]), .O(n32));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut.LUT_INIT = 16'h8421;
    SB_LUT4 i4335_3_lut (.I0(\REG.mem_47_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n18), .I3(GND_net), .O(n5718));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4336_3_lut (.I0(\REG.mem_47_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n18), .I3(GND_net), .O(n5719));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n4335), 
            .I3(debug_led3), .O(n10406));   // src/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i1_3_lut (.I0(is_fifo_empty_flag), .I1(fifo_write_cmd), .I2(n32), 
            .I3(GND_net), .O(n24));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i9060_4_lut (.I0(rd_addr_p1_w_adj_123[2]), .I1(n14025), .I2(wr_addr_r_adj_118[2]), 
            .I3(wr_addr_r_adj_118[1]), .O(n10897));
    defparam i9060_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_86 (.I0(reset_all_w), .I1(n10897), .I2(n24), 
            .I3(n4_adj_58), .O(n10786));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_adj_86.LUT_INIT = 16'hfbfa;
    SB_LUT4 i4337_3_lut (.I0(\REG.mem_47_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n18), .I3(GND_net), .O(n5720));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4662_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[1]), .I2(GND_net), 
            .I3(GND_net), .O(n6045));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4662_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4338_3_lut (.I0(\REG.mem_48_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n17), .I3(GND_net), .O(n5721));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4339_3_lut (.I0(\REG.mem_48_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n17), .I3(GND_net), .O(n5722));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4340_3_lut (.I0(\REG.mem_48_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n17), .I3(GND_net), .O(n5723));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4341_3_lut (.I0(\REG.mem_48_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n17), .I3(GND_net), .O(n5724));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4342_3_lut (.I0(\REG.mem_48_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n17), .I3(GND_net), .O(n5725));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4343_3_lut (.I0(\REG.mem_48_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n17), .I3(GND_net), .O(n5726));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4344_3_lut (.I0(\REG.mem_48_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n17), .I3(GND_net), .O(n5727));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4345_3_lut (.I0(\REG.mem_48_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n17), .I3(GND_net), .O(n5728));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4346_3_lut (.I0(\REG.mem_48_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n17), .I3(GND_net), .O(n5729));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4347_3_lut (.I0(\REG.mem_48_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n17), .I3(GND_net), .O(n5730));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4671_3_lut (.I0(rx_buf_byte[7]), .I1(rx_shift_reg[7]), .I2(n3495), 
            .I3(GND_net), .O(n6054));   // src/spi.v(76[8] 221[4])
    defparam i4671_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4672_3_lut (.I0(rx_buf_byte[6]), .I1(rx_shift_reg[6]), .I2(n3495), 
            .I3(GND_net), .O(n6055));   // src/spi.v(76[8] 221[4])
    defparam i4672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4246_3_lut (.I0(\REG.mem_42_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n23), .I3(GND_net), .O(n5629));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4348_3_lut (.I0(\REG.mem_48_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n17), .I3(GND_net), .O(n5731));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1186_1260_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_65), .I3(n10174), .O(n127)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4247_3_lut (.I0(\REG.mem_42_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n23), .I3(GND_net), .O(n5630));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4248_3_lut (.I0(\REG.mem_42_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n23), .I3(GND_net), .O(n5631));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4349_3_lut (.I0(\REG.mem_48_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n17), .I3(GND_net), .O(n5732));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4249_3_lut (.I0(\REG.mem_42_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n23), .I3(GND_net), .O(n5632));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4673_3_lut (.I0(rx_buf_byte[5]), .I1(rx_shift_reg[5]), .I2(n3495), 
            .I3(GND_net), .O(n6056));   // src/spi.v(76[8] 221[4])
    defparam i4673_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4350_3_lut (.I0(\REG.mem_48_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n17), .I3(GND_net), .O(n5733));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4250_3_lut (.I0(\REG.mem_42_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n23), .I3(GND_net), .O(n5633));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4351_3_lut (.I0(\REG.mem_48_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n17), .I3(GND_net), .O(n5734));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4352_3_lut (.I0(\REG.mem_48_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n17), .I3(GND_net), .O(n5735));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4674_3_lut (.I0(rx_buf_byte[4]), .I1(rx_shift_reg[4]), .I2(n3495), 
            .I3(GND_net), .O(n6057));   // src/spi.v(76[8] 221[4])
    defparam i4674_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4675_3_lut (.I0(rx_buf_byte[3]), .I1(rx_shift_reg[3]), .I2(n3495), 
            .I3(GND_net), .O(n6058));   // src/spi.v(76[8] 221[4])
    defparam i4675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4676_3_lut (.I0(rx_buf_byte[2]), .I1(rx_shift_reg[2]), .I2(n3495), 
            .I3(GND_net), .O(n6059));   // src/spi.v(76[8] 221[4])
    defparam i4676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4251_3_lut (.I0(\REG.mem_42_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n23), .I3(GND_net), .O(n5634));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4353_3_lut (.I0(\REG.mem_48_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n17), .I3(GND_net), .O(n5736));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4252_3_lut (.I0(\REG.mem_42_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n23), .I3(GND_net), .O(n5635));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4253_3_lut (.I0(\REG.mem_42_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n23), .I3(GND_net), .O(n5636));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4677_3_lut (.I0(rx_buf_byte[1]), .I1(rx_shift_reg[1]), .I2(n3495), 
            .I3(GND_net), .O(n6060));   // src/spi.v(76[8] 221[4])
    defparam i4677_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 reset_all_w_I_0_1_lut (.I0(reset_all_w), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(RESET_c));   // src/top.v(295[16:28])
    defparam reset_all_w_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4254_3_lut (.I0(\REG.mem_42_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n23), .I3(GND_net), .O(n5637));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4255_3_lut (.I0(\REG.mem_43_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n22), .I3(GND_net), .O(n5638));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4256_3_lut (.I0(\REG.mem_43_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n22), .I3(GND_net), .O(n5639));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4257_3_lut (.I0(\REG.mem_43_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n22), .I3(GND_net), .O(n5640));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4258_3_lut (.I0(\REG.mem_43_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n22), .I3(GND_net), .O(n5641));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4691_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[1]), .I2(n4_adj_77), 
            .I3(n4253), .O(n6074));   // src/uart_rx.v(49[10] 144[8])
    defparam i4691_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4692_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[2]), .I2(n4), 
            .I3(n4248), .O(n6075));   // src/uart_rx.v(49[10] 144[8])
    defparam i4692_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1655_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n3022));   // src/top.v(1074[8] 1141[4])
    defparam i1655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4259_3_lut (.I0(\REG.mem_43_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n22), .I3(GND_net), .O(n5642));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4694_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[3]), .I2(n4), 
            .I3(n4253), .O(n6077));   // src/uart_rx.v(49[10] 144[8])
    defparam i4694_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4695_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[4]), .I2(n4_adj_78), 
            .I3(n4248), .O(n6078));   // src/uart_rx.v(49[10] 144[8])
    defparam i4695_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4696_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[5]), .I2(n4_adj_78), 
            .I3(n4253), .O(n6079));   // src/uart_rx.v(49[10] 144[8])
    defparam i4696_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4260_3_lut (.I0(\REG.mem_43_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n22), .I3(GND_net), .O(n5643));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4260_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF start_tx_81 (.Q(r_SM_Main_2__N_844[0]), .C(SLM_CLK_c), .D(n6106));   // src/top.v(910[8] 928[4])
    SB_LUT4 i4698_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[6]), .I2(n7473), 
            .I3(n4248), .O(n6081));   // src/uart_rx.v(49[10] 144[8])
    defparam i4698_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i4699_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[7]), .I2(n7473), 
            .I3(n4253), .O(n6082));   // src/uart_rx.v(49[10] 144[8])
    defparam i4699_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i4705_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[0]), .I2(\mem_LUT.data_raw_r [0]), 
            .I3(n4459), .O(n6088));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4705_4_lut.LUT_INIT = 16'h5044;
    SB_CARRY led_counter_1186_1260_add_4_5 (.CI(n10174), .I0(GND_net), .I1(n22_adj_65), 
            .CO(n10175));
    SB_LUT4 i4261_3_lut (.I0(\REG.mem_43_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n22), .I3(GND_net), .O(n5644));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_87 (.I0(buffer_switch_done_latched), .I1(n843), 
            .I2(n771), .I3(GND_net), .O(n10277));
    defparam i1_3_lut_adj_87.LUT_INIT = 16'heaea;
    SB_LUT4 i4262_3_lut (.I0(\REG.mem_43_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n22), .I3(GND_net), .O(n5645));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4370_3_lut (.I0(\REG.mem_50_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n15_adj_60), .I3(GND_net), .O(n5753));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4263_3_lut (.I0(\REG.mem_43_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n22), .I3(GND_net), .O(n5646));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4264_3_lut (.I0(\REG.mem_43_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n22), .I3(GND_net), .O(n5647));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4265_3_lut (.I0(\REG.mem_43_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n22), .I3(GND_net), .O(n5648));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4266_3_lut (.I0(\REG.mem_43_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n22), .I3(GND_net), .O(n5649));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4267_3_lut (.I0(\REG.mem_43_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n22), .I3(GND_net), .O(n5650));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4268_3_lut (.I0(\REG.mem_43_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n22), .I3(GND_net), .O(n5651));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4268_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF spi_start_transfer_r_84 (.Q(spi_start_transfer_r), .C(SLM_CLK_c), 
           .D(n3022));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 i3504_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[3]), .I2(\mem_LUT.data_raw_r [3]), 
            .I3(n4459), .O(n4887));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i3504_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4269_3_lut (.I0(\REG.mem_43_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n22), .I3(GND_net), .O(n5652));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4374_3_lut (.I0(\REG.mem_50_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n15_adj_60), .I3(GND_net), .O(n5757));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4375_3_lut (.I0(\REG.mem_50_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n15_adj_60), .I3(GND_net), .O(n5758));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4376_3_lut (.I0(\REG.mem_50_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n15_adj_60), .I3(GND_net), .O(n5759));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4377_3_lut (.I0(\REG.mem_50_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n15_adj_60), .I3(GND_net), .O(n5760));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4378_3_lut (.I0(\REG.mem_50_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n15_adj_60), .I3(GND_net), .O(n5761));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4722_3_lut (.I0(pc_data_rx[0]), .I1(r_Rx_Data), .I2(n10345), 
            .I3(GND_net), .O(n6105));   // src/uart_rx.v(49[10] 144[8])
    defparam i4722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4270_3_lut (.I0(\REG.mem_43_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n22), .I3(GND_net), .O(n5653));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4379_3_lut (.I0(\REG.mem_50_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n15_adj_60), .I3(GND_net), .O(n5762));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4271_3_lut (.I0(\REG.mem_44_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n21), .I3(GND_net), .O(n5654));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10377_2_lut (.I0(is_fifo_empty_flag), .I1(tx_uart_active_flag), 
            .I2(GND_net), .I3(GND_net), .O(start_tx_N_64));
    defparam i10377_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i4380_3_lut (.I0(\REG.mem_50_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n15_adj_60), .I3(GND_net), .O(n5763));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4272_3_lut (.I0(\REG.mem_44_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n21), .I3(GND_net), .O(n5655));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4381_3_lut (.I0(\REG.mem_50_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n15_adj_60), .I3(GND_net), .O(n5764));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4381_3_lut.LUT_INIT = 16'hcaca;
    GND i1 (.Y(GND_net));
    SB_LUT4 i4273_3_lut (.I0(\REG.mem_44_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n21), .I3(GND_net), .O(n5656));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4382_3_lut (.I0(\REG.mem_50_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n15_adj_60), .I3(GND_net), .O(n5765));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4383_3_lut (.I0(\REG.mem_50_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n15_adj_60), .I3(GND_net), .O(n5766));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9080_4_lut (.I0(n1), .I1(fifo_read_cmd), .I2(wr_addr_r_adj_118[1]), 
            .I3(rd_addr_r_adj_121[1]), .O(n10917));
    defparam i9080_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i4384_3_lut (.I0(\REG.mem_50_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n15_adj_60), .I3(GND_net), .O(n5767));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4274_3_lut (.I0(\REG.mem_44_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n21), .I3(GND_net), .O(n5657));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4274_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4385_3_lut (.I0(\REG.mem_50_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n15_adj_60), .I3(GND_net), .O(n5768));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4275_3_lut (.I0(\REG.mem_44_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n21), .I3(GND_net), .O(n5658));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_88 (.I0(reset_all_w), .I1(n15), .I2(wr_fifo_en_w), 
            .I3(n10226), .O(n10430));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_adj_88.LUT_INIT = 16'h5444;
    SB_LUT4 i4276_3_lut (.I0(\REG.mem_44_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n21), .I3(GND_net), .O(n5659));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4386_3_lut (.I0(\REG.mem_50_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n15_adj_60), .I3(GND_net), .O(n5769));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4277_3_lut (.I0(\REG.mem_44_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n21), .I3(GND_net), .O(n5660));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4387_3_lut (.I0(\REG.mem_50_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n15_adj_60), .I3(GND_net), .O(n5770));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut (.I0(tx_shift_reg[0]), .I1(n2086), .I2(n4319), .I3(tx_data_byte[0]), 
            .O(n10428));   // src/spi.v(76[8] 221[4])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i4388_3_lut (.I0(\REG.mem_50_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n15_adj_60), .I3(GND_net), .O(n5771));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9035_2_lut (.I0(n63), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n10871));
    defparam i9035_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 led_counter_1186_1260_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_64), .I3(n10173), .O(n128)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19_4_lut (.I0(n4245), .I1(n12063), .I2(state[3]), .I3(n10871), 
            .O(n10514));   // src/timing_controller.v(56[8] 132[4])
    defparam i19_4_lut.LUT_INIT = 16'hfcac;
    SB_DFF tx_data_byte_r_i0_i5 (.Q(tx_data_byte[5]), .C(SLM_CLK_c), .D(n5970));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 i4744_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[1]), .I2(\mem_LUT.data_raw_r [1]), 
            .I3(n4459), .O(n6127));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4744_4_lut.LUT_INIT = 16'h5044;
    SB_CARRY led_counter_1186_1260_add_4_4 (.CI(n10173), .I0(GND_net), .I1(n23_adj_64), 
            .CO(n10174));
    SB_LUT4 led_counter_1186_1260_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_63), .I3(n10172), .O(n129)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_3 (.CI(n10172), .I0(GND_net), .I1(n24_adj_63), 
            .CO(n10173));
    SB_LUT4 led_counter_1186_1260_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_62), .I3(VCC_net), .O(n130)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(n25_adj_62), .CO(n10172));
    SB_LUT4 led_counter_1186_1260_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(DEBUG_0_c_24), .I3(n10195), .O(n106)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 led_counter_1186_1260_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n2_adj_75), .I3(n10194), .O(n107)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_25 (.CI(n10194), .I0(GND_net), 
            .I1(n2_adj_75), .CO(n10195));
    SB_LUT4 led_counter_1186_1260_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3), .I3(n10193), .O(n108)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_24 (.CI(n10193), .I0(GND_net), 
            .I1(n3), .CO(n10194));
    SB_LUT4 led_counter_1186_1260_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_74), .I3(n10192), .O(n109)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_23 (.CI(n10192), .I0(GND_net), 
            .I1(n4_adj_74), .CO(n10193));
    SB_LUT4 led_counter_1186_1260_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5), .I3(n10191), .O(n110)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_22 (.CI(n10191), .I0(GND_net), 
            .I1(n5), .CO(n10192));
    SB_LUT4 led_counter_1186_1260_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6), .I3(n10190), .O(n111)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_21 (.CI(n10190), .I0(GND_net), 
            .I1(n6), .CO(n10191));
    SB_LUT4 led_counter_1186_1260_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7), .I3(n10189), .O(n112)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_20 (.CI(n10189), .I0(GND_net), 
            .I1(n7), .CO(n10190));
    SB_LUT4 led_counter_1186_1260_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_73), .I3(n10188), .O(n113)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_19 (.CI(n10188), .I0(GND_net), 
            .I1(n8_adj_73), .CO(n10189));
    SB_LUT4 led_counter_1186_1260_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9), .I3(n10187), .O(n114)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_18 (.CI(n10187), .I0(GND_net), 
            .I1(n9), .CO(n10188));
    SB_LUT4 led_counter_1186_1260_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_72), .I3(n10186), .O(n115)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_17 (.CI(n10186), .I0(GND_net), 
            .I1(n10_adj_72), .CO(n10187));
    SB_LUT4 led_counter_1186_1260_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11), .I3(n10185), .O(n116)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_16 (.CI(n10185), .I0(GND_net), 
            .I1(n11), .CO(n10186));
    SB_LUT4 led_counter_1186_1260_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12), .I3(n10184), .O(n117)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_15 (.CI(n10184), .I0(GND_net), 
            .I1(n12), .CO(n10185));
    SB_LUT4 i1_3_lut_adj_89 (.I0(reset_clk_counter[3]), .I1(reset_clk_counter[2]), 
            .I2(n10064), .I3(GND_net), .O(n10293));
    defparam i1_3_lut_adj_89.LUT_INIT = 16'ha9a9;
    SB_LUT4 led_counter_1186_1260_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13), .I3(n10183), .O(n118)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_14 (.CI(n10183), .I0(GND_net), 
            .I1(n13), .CO(n10184));
    SB_LUT4 led_counter_1186_1260_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14), .I3(n10182), .O(n119)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_IO FIFO_D1_pad (.PACKAGE_PIN(FIFO_D1), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D1_c_1));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D1_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D1_pad.PULLUP = 1'b0;
    defparam FIFO_D1_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D2_pad (.PACKAGE_PIN(FIFO_D2), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D2_c_2));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D2_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D2_pad.PULLUP = 1'b0;
    defparam FIFO_D2_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D3_pad (.PACKAGE_PIN(FIFO_D3), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D3_c_3));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D3_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D3_pad.PULLUP = 1'b0;
    defparam FIFO_D3_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY led_counter_1186_1260_add_4_13 (.CI(n10182), .I0(GND_net), 
            .I1(n14), .CO(n10183));
    SB_IO FIFO_D4_pad (.PACKAGE_PIN(FIFO_D4), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D4_c_4));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D4_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D4_pad.PULLUP = 1'b0;
    defparam FIFO_D4_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D5_pad (.PACKAGE_PIN(FIFO_D5), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D5_c_5));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D5_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D5_pad.PULLUP = 1'b0;
    defparam FIFO_D5_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D6_pad (.PACKAGE_PIN(FIFO_D6), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D6_c_6));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D6_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D6_pad.PULLUP = 1'b0;
    defparam FIFO_D6_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D7_pad (.PACKAGE_PIN(FIFO_D7), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D7_c_7));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D7_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D7_pad.PULLUP = 1'b0;
    defparam FIFO_D7_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D8_pad (.PACKAGE_PIN(FIFO_D8), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D8_c_8));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D8_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D8_pad.PULLUP = 1'b0;
    defparam FIFO_D8_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D9_pad (.PACKAGE_PIN(FIFO_D9), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D9_c_9));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D9_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D9_pad.PULLUP = 1'b0;
    defparam FIFO_D9_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D10_pad (.PACKAGE_PIN(FIFO_D10), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D10_c_10));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D10_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D10_pad.PULLUP = 1'b0;
    defparam FIFO_D10_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D11_pad (.PACKAGE_PIN(FIFO_D11), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D11_c_11));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D11_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D11_pad.PULLUP = 1'b0;
    defparam FIFO_D11_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D12_pad (.PACKAGE_PIN(FIFO_D12), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D12_c_12));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D12_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D12_pad.PULLUP = 1'b0;
    defparam FIFO_D12_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D13_pad (.PACKAGE_PIN(FIFO_D13), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D13_c_13));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D13_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D13_pad.PULLUP = 1'b0;
    defparam FIFO_D13_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D14_pad (.PACKAGE_PIN(FIFO_D14), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D14_c_14));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D14_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D14_pad.PULLUP = 1'b0;
    defparam FIFO_D14_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D15_pad (.PACKAGE_PIN(FIFO_D15), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D15_c_15));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D15_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D15_pad.PULLUP = 1'b0;
    defparam FIFO_D15_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D15_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO FIFO_CLK_pad (.PACKAGE_PIN(FIFO_CLK), .OUTPUT_ENABLE(VCC_net), 
            .GLOBAL_BUFFER_OUTPUT(FIFO_CLK_c));   // src/top.v(84[12:20])
    defparam FIFO_CLK_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_CLK_pad.PULLUP = 1'b0;
    defparam FIFO_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_1_c_pad (.PACKAGE_PIN(FR_RXF), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(DEBUG_1_c_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_1_c_pad.PIN_TYPE = 6'b000001;
    defparam DEBUG_1_c_pad.PULLUP = 1'b0;
    defparam DEBUG_1_c_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_1_c_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SOUT_pad (.PACKAGE_PIN(SOUT), .OUTPUT_ENABLE(VCC_net), .D_IN_0(SOUT_c)) /* synthesis IO_FF_IN=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SOUT_pad.PIN_TYPE = 6'b000001;
    defparam SOUT_pad.PULLUP = 1'b0;
    defparam SOUT_pad.NEG_TRIGGER = 1'b0;
    defparam SOUT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UART_RX_pad (.PACKAGE_PIN(UART_RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(UART_RX_c)) /* synthesis IO_FF_IN=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UART_RX_pad.PIN_TYPE = 6'b000001;
    defparam UART_RX_pad.PULLUP = 1'b0;
    defparam UART_RX_pad.NEG_TRIGGER = 1'b0;
    defparam UART_RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_SYSCLK_pad (.PACKAGE_PIN(ICE_SYSCLK), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ICE_SYSCLK_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_SYSCLK_pad.PIN_TYPE = 6'b000001;
    defparam ICE_SYSCLK_pad.PULLUP = 1'b0;
    defparam ICE_SYSCLK_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_SYSCLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CREST_pad (.PACKAGE_PIN(ICE_CREST), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CREST_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CREST_pad.PULLUP = 1'b0;
    defparam ICE_CREST_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CREST_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CDONE_pad (.PACKAGE_PIN(ICE_CDONE), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CDONE_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CDONE_pad.PULLUP = 1'b0;
    defparam ICE_CDONE_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CDONE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CLK_pad (.PACKAGE_PIN(ICE_CLK), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CLK_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CLK_pad.PULLUP = 1'b0;
    defparam ICE_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_9_pad (.PACKAGE_PIN(DEBUG_9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_9_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_9_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_9_pad.PULLUP = 1'b0;
    defparam DEBUG_9_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_8_pad (.PACKAGE_PIN(DEBUG_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_8_c_0_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_8_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_8_pad.PULLUP = 1'b0;
    defparam DEBUG_8_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_6_pad (.PACKAGE_PIN(DEBUG_6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_6_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_6_pad.PULLUP = 1'b0;
    defparam DEBUG_6_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_5_pad (.PACKAGE_PIN(DEBUG_5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_5_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_5_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_5_pad.PULLUP = 1'b0;
    defparam DEBUG_5_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_3_pad (.PACKAGE_PIN(DEBUG_3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_3_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_3_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_3_pad.PULLUP = 1'b0;
    defparam DEBUG_3_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_2_pad (.PACKAGE_PIN(DEBUG_2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_2_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_2_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_2_pad.PULLUP = 1'b0;
    defparam DEBUG_2_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_1_pad (.PACKAGE_PIN(DEBUG_1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_1_c_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_1_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_1_pad.PULLUP = 1'b0;
    defparam DEBUG_1_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_0_pad (.PACKAGE_PIN(DEBUG_0), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_0_c_24));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_0_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_0_pad.PULLUP = 1'b0;
    defparam DEBUG_0_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_SIWU_pad (.PACKAGE_PIN(FT_SIWU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_SIWU_pad.PIN_TYPE = 6'b011001;
    defparam FT_SIWU_pad.PULLUP = 1'b0;
    defparam FT_SIWU_pad.NEG_TRIGGER = 1'b0;
    defparam FT_SIWU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_WR_pad (.PACKAGE_PIN(FT_WR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_WR_pad.PIN_TYPE = 6'b011001;
    defparam FT_WR_pad.PULLUP = 1'b0;
    defparam FT_WR_pad.NEG_TRIGGER = 1'b0;
    defparam FT_WR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_RD_pad (.PACKAGE_PIN(FT_RD), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_2_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_RD_pad.PIN_TYPE = 6'b011001;
    defparam FT_RD_pad.PULLUP = 1'b0;
    defparam FT_RD_pad.NEG_TRIGGER = 1'b0;
    defparam FT_RD_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_OE_pad (.PACKAGE_PIN(FT_OE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(FT_OE_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_OE_pad.PIN_TYPE = 6'b011001;
    defparam FT_OE_pad.PULLUP = 1'b0;
    defparam FT_OE_pad.NEG_TRIGGER = 1'b0;
    defparam FT_OE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA10_pad (.PACKAGE_PIN(DATA10), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA10_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA10_pad.PIN_TYPE = 6'b011001;
    defparam DATA10_pad.PULLUP = 1'b0;
    defparam DATA10_pad.NEG_TRIGGER = 1'b0;
    defparam DATA10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA9_pad (.PACKAGE_PIN(DATA9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA9_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA9_pad.PIN_TYPE = 6'b011001;
    defparam DATA9_pad.PULLUP = 1'b0;
    defparam DATA9_pad.NEG_TRIGGER = 1'b0;
    defparam DATA9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA11_pad (.PACKAGE_PIN(DATA11), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA11_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA11_pad.PIN_TYPE = 6'b011001;
    defparam DATA11_pad.PULLUP = 1'b0;
    defparam DATA11_pad.NEG_TRIGGER = 1'b0;
    defparam DATA11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA12_pad (.PACKAGE_PIN(DATA12), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA12_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA12_pad.PIN_TYPE = 6'b011001;
    defparam DATA12_pad.PULLUP = 1'b0;
    defparam DATA12_pad.NEG_TRIGGER = 1'b0;
    defparam DATA12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA13_pad (.PACKAGE_PIN(DATA13), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA13_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA13_pad.PIN_TYPE = 6'b011001;
    defparam DATA13_pad.PULLUP = 1'b0;
    defparam DATA13_pad.NEG_TRIGGER = 1'b0;
    defparam DATA13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA14_pad (.PACKAGE_PIN(DATA14), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA14_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA14_pad.PIN_TYPE = 6'b011001;
    defparam DATA14_pad.PULLUP = 1'b0;
    defparam DATA14_pad.NEG_TRIGGER = 1'b0;
    defparam DATA14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA8_pad (.PACKAGE_PIN(DATA8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA8_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA8_pad.PIN_TYPE = 6'b011001;
    defparam DATA8_pad.PULLUP = 1'b0;
    defparam DATA8_pad.NEG_TRIGGER = 1'b0;
    defparam DATA8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA15_pad (.PACKAGE_PIN(DATA15), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA15_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA15_pad.PIN_TYPE = 6'b011001;
    defparam DATA15_pad.PULLUP = 1'b0;
    defparam DATA15_pad.NEG_TRIGGER = 1'b0;
    defparam DATA15_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA16_pad (.PACKAGE_PIN(DATA16), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA16_pad.PIN_TYPE = 6'b011001;
    defparam DATA16_pad.PULLUP = 1'b0;
    defparam DATA16_pad.NEG_TRIGGER = 1'b0;
    defparam DATA16_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA7_pad (.PACKAGE_PIN(DATA7), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA7_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA7_pad.PIN_TYPE = 6'b011001;
    defparam DATA7_pad.PULLUP = 1'b0;
    defparam DATA7_pad.NEG_TRIGGER = 1'b0;
    defparam DATA7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA17_pad (.PACKAGE_PIN(DATA17), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA17_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA17_pad.PIN_TYPE = 6'b011001;
    defparam DATA17_pad.PULLUP = 1'b0;
    defparam DATA17_pad.NEG_TRIGGER = 1'b0;
    defparam DATA17_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA18_pad (.PACKAGE_PIN(DATA18), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA18_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA18_pad.PIN_TYPE = 6'b011001;
    defparam DATA18_pad.PULLUP = 1'b0;
    defparam DATA18_pad.NEG_TRIGGER = 1'b0;
    defparam DATA18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA6_pad (.PACKAGE_PIN(DATA6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA6_pad.PIN_TYPE = 6'b011001;
    defparam DATA6_pad.PULLUP = 1'b0;
    defparam DATA6_pad.NEG_TRIGGER = 1'b0;
    defparam DATA6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA19_pad (.PACKAGE_PIN(DATA19), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA19_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA19_pad.PIN_TYPE = 6'b011001;
    defparam DATA19_pad.PULLUP = 1'b0;
    defparam DATA19_pad.NEG_TRIGGER = 1'b0;
    defparam DATA19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA20_pad (.PACKAGE_PIN(DATA20), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA20_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA20_pad.PIN_TYPE = 6'b011001;
    defparam DATA20_pad.PULLUP = 1'b0;
    defparam DATA20_pad.NEG_TRIGGER = 1'b0;
    defparam DATA20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA5_pad (.PACKAGE_PIN(DATA5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA5_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA5_pad.PIN_TYPE = 6'b011001;
    defparam DATA5_pad.PULLUP = 1'b0;
    defparam DATA5_pad.NEG_TRIGGER = 1'b0;
    defparam DATA5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA21_pad (.PACKAGE_PIN(DATA21), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA5_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA21_pad.PIN_TYPE = 6'b011001;
    defparam DATA21_pad.PULLUP = 1'b0;
    defparam DATA21_pad.NEG_TRIGGER = 1'b0;
    defparam DATA21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA22_pad (.PACKAGE_PIN(DATA22), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA22_pad.PIN_TYPE = 6'b011001;
    defparam DATA22_pad.PULLUP = 1'b0;
    defparam DATA22_pad.NEG_TRIGGER = 1'b0;
    defparam DATA22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA4_pad (.PACKAGE_PIN(DATA4), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA20_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA4_pad.PIN_TYPE = 6'b011001;
    defparam DATA4_pad.PULLUP = 1'b0;
    defparam DATA4_pad.NEG_TRIGGER = 1'b0;
    defparam DATA4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA23_pad (.PACKAGE_PIN(DATA23), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA7_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA23_pad.PIN_TYPE = 6'b011001;
    defparam DATA23_pad.PULLUP = 1'b0;
    defparam DATA23_pad.NEG_TRIGGER = 1'b0;
    defparam DATA23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA24_pad (.PACKAGE_PIN(DATA24), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA8_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA24_pad.PIN_TYPE = 6'b011001;
    defparam DATA24_pad.PULLUP = 1'b0;
    defparam DATA24_pad.NEG_TRIGGER = 1'b0;
    defparam DATA24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA3_pad (.PACKAGE_PIN(DATA3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA19_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA3_pad.PIN_TYPE = 6'b011001;
    defparam DATA3_pad.PULLUP = 1'b0;
    defparam DATA3_pad.NEG_TRIGGER = 1'b0;
    defparam DATA3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 led_counter_1186_1260_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_71), .I3(n10181), .O(n120)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_IO DATA25_pad (.PACKAGE_PIN(DATA25), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA9_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA25_pad.PIN_TYPE = 6'b011001;
    defparam DATA25_pad.PULLUP = 1'b0;
    defparam DATA25_pad.NEG_TRIGGER = 1'b0;
    defparam DATA25_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA26_pad (.PACKAGE_PIN(DATA26), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA10_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA26_pad.PIN_TYPE = 6'b011001;
    defparam DATA26_pad.PULLUP = 1'b0;
    defparam DATA26_pad.NEG_TRIGGER = 1'b0;
    defparam DATA26_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA2_pad (.PACKAGE_PIN(DATA2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA18_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA2_pad.PIN_TYPE = 6'b011001;
    defparam DATA2_pad.PULLUP = 1'b0;
    defparam DATA2_pad.NEG_TRIGGER = 1'b0;
    defparam DATA2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA27_pad (.PACKAGE_PIN(DATA27), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA11_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA27_pad.PIN_TYPE = 6'b011001;
    defparam DATA27_pad.PULLUP = 1'b0;
    defparam DATA27_pad.NEG_TRIGGER = 1'b0;
    defparam DATA27_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA28_pad (.PACKAGE_PIN(DATA28), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA12_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA28_pad.PIN_TYPE = 6'b011001;
    defparam DATA28_pad.PULLUP = 1'b0;
    defparam DATA28_pad.NEG_TRIGGER = 1'b0;
    defparam DATA28_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA1_pad (.PACKAGE_PIN(DATA1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA17_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA1_pad.PIN_TYPE = 6'b011001;
    defparam DATA1_pad.PULLUP = 1'b0;
    defparam DATA1_pad.NEG_TRIGGER = 1'b0;
    defparam DATA1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA29_pad (.PACKAGE_PIN(DATA29), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA13_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA29_pad.PIN_TYPE = 6'b011001;
    defparam DATA29_pad.PULLUP = 1'b0;
    defparam DATA29_pad.NEG_TRIGGER = 1'b0;
    defparam DATA29_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA30_pad (.PACKAGE_PIN(DATA30), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA14_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA30_pad.PIN_TYPE = 6'b011001;
    defparam DATA30_pad.PULLUP = 1'b0;
    defparam DATA30_pad.NEG_TRIGGER = 1'b0;
    defparam DATA30_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA0_pad (.PACKAGE_PIN(DATA0), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA0_pad.PIN_TYPE = 6'b011001;
    defparam DATA0_pad.PULLUP = 1'b0;
    defparam DATA0_pad.NEG_TRIGGER = 1'b0;
    defparam DATA0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY led_counter_1186_1260_add_4_12 (.CI(n10181), .I0(GND_net), 
            .I1(n15_adj_71), .CO(n10182));
    SB_IO DATA31_pad (.PACKAGE_PIN(DATA31), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA15_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA31_pad.PIN_TYPE = 6'b011001;
    defparam DATA31_pad.PULLUP = 1'b0;
    defparam DATA31_pad.NEG_TRIGGER = 1'b0;
    defparam DATA31_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO VALID_pad (.PACKAGE_PIN(VALID), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_9_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam VALID_pad.PIN_TYPE = 6'b011001;
    defparam VALID_pad.PULLUP = 1'b0;
    defparam VALID_pad.NEG_TRIGGER = 1'b0;
    defparam VALID_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SYNC_pad (.PACKAGE_PIN(SYNC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SYNC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SYNC_pad.PIN_TYPE = 6'b011001;
    defparam SYNC_pad.PULLUP = 1'b0;
    defparam SYNC_pad.NEG_TRIGGER = 1'b0;
    defparam SYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INVERT_pad (.PACKAGE_PIN(INVERT), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INVERT_c_3)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INVERT_pad.PIN_TYPE = 6'b011001;
    defparam INVERT_pad.PULLUP = 1'b0;
    defparam INVERT_pad.NEG_TRIGGER = 1'b0;
    defparam INVERT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SLM_CLK_pad (.PACKAGE_PIN(SLM_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SLM_CLK_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SLM_CLK_pad.PIN_TYPE = 6'b011001;
    defparam SLM_CLK_pad.PULLUP = 1'b0;
    defparam SLM_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam SLM_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO RESET_pad (.PACKAGE_PIN(RESET), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(RESET_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RESET_pad.PIN_TYPE = 6'b011001;
    defparam RESET_pad.PULLUP = 1'b0;
    defparam RESET_pad.NEG_TRIGGER = 1'b0;
    defparam RESET_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UPDATE_pad (.PACKAGE_PIN(UPDATE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(UPDATE_c_2));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UPDATE_pad.PIN_TYPE = 6'b011001;
    defparam UPDATE_pad.PULLUP = 1'b0;
    defparam UPDATE_pad.NEG_TRIGGER = 1'b0;
    defparam UPDATE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SDAT_pad (.PACKAGE_PIN(SDAT), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SDAT_c_15)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SDAT_pad.PIN_TYPE = 6'b011001;
    defparam SDAT_pad.PULLUP = 1'b0;
    defparam SDAT_pad.NEG_TRIGGER = 1'b0;
    defparam SDAT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SCK_pad (.PACKAGE_PIN(SCK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SCK_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SCK_pad.PIN_TYPE = 6'b011001;
    defparam SCK_pad.PULLUP = 1'b0;
    defparam SCK_pad.NEG_TRIGGER = 1'b0;
    defparam SCK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SEN_pad (.PACKAGE_PIN(SEN), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SEN_c_1)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SEN_pad.PIN_TYPE = 6'b011001;
    defparam SEN_pad.PULLUP = 1'b0;
    defparam SEN_pad.NEG_TRIGGER = 1'b0;
    defparam SEN_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UART_TX_pad (.PACKAGE_PIN(UART_TX), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(UART_TX_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UART_TX_pad.PIN_TYPE = 6'b011001;
    defparam UART_TX_pad.PULLUP = 1'b0;
    defparam UART_TX_pad.NEG_TRIGGER = 1'b0;
    defparam UART_TX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i3556_2_lut (.I0(is_tx_fifo_full_flag), .I1(spi_rx_byte_ready), 
            .I2(GND_net), .I3(GND_net), .O(n4939));   // src/top.v(889[8] 898[4])
    defparam i3556_2_lut.LUT_INIT = 16'h4444;
    SB_DFF tx_addr_byte_r_i0_i0 (.Q(tx_addr_byte[0]), .C(SLM_CLK_c), .D(n4923));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 led_counter_1186_1260_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16), .I3(n10180), .O(n121)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_11 (.CI(n10180), .I0(GND_net), 
            .I1(n16), .CO(n10181));
    SB_LUT4 led_counter_1186_1260_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_70), .I3(n10179), .O(n122)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_10 (.CI(n10179), .I0(GND_net), 
            .I1(n17_adj_70), .CO(n10180));
    SB_DFF uart_rx_complete_rising_edge_82 (.Q(uart_rx_complete_rising_edge), 
           .C(SLM_CLK_c), .D(n4909));   // src/top.v(1065[8] 1071[4])
    SB_LUT4 led_counter_1186_1260_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_69), .I3(n10178), .O(n123)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF tx_addr_byte_r_i0_i1 (.Q(tx_addr_byte[1]), .C(SLM_CLK_c), .D(n5533));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_addr_byte_r_i0_i2 (.Q(tx_addr_byte[2]), .C(SLM_CLK_c), .D(n5532));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_addr_byte_r_i0_i3 (.Q(tx_addr_byte[3]), .C(SLM_CLK_c), .D(n5531));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_addr_byte_r_i0_i4 (.Q(tx_addr_byte[4]), .C(SLM_CLK_c), .D(n5530));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_addr_byte_r_i0_i5 (.Q(tx_addr_byte[5]), .C(SLM_CLK_c), .D(n5529));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_addr_byte_r_i0_i6 (.Q(tx_addr_byte[6]), .C(SLM_CLK_c), .D(n5528));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_addr_byte_r_i0_i7 (.Q(tx_addr_byte[7]), .C(SLM_CLK_c), .D(n5527));   // src/top.v(1074[8] 1141[4])
    SB_CARRY led_counter_1186_1260_add_4_9 (.CI(n10178), .I0(GND_net), .I1(n18_adj_69), 
            .CO(n10179));
    SB_DFF tx_data_byte_r_i0_i6 (.Q(tx_data_byte[6]), .C(SLM_CLK_c), .D(n5510));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 i3559_3_lut (.I0(tx_data_byte[7]), .I1(pc_data_rx[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4942));   // src/top.v(1074[8] 1141[4])
    defparam i3559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4453_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[6]), .I2(GND_net), 
            .I3(GND_net), .O(n5836));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4453_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4454_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5837));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4454_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4455_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5838));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4455_2_lut.LUT_INIT = 16'h4444;
    SB_DFF reset_clk_counter_i3_1187__i0 (.Q(reset_clk_counter[0]), .C(SLM_CLK_c), 
           .D(n25_adj_76));   // src/top.v(259[27:51])
    SB_LUT4 i4456_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5839));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4456_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3499_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[2]), .I2(\mem_LUT.data_raw_r [2]), 
            .I3(n4459), .O(n4882));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i3499_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4458_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5841));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4458_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i954_4_lut (.I0(n2034), .I1(n7568), .I2(state[3]), .I3(n63), 
            .O(n1879));   // src/timing_controller.v(51[11:16])
    defparam i954_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i4459_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5842));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4459_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3181_4_lut (.I0(n63), .I1(n4192), .I2(n7568), .I3(state[3]), 
            .O(n1774));   // src/timing_controller.v(51[11:16])
    defparam i3181_4_lut.LUT_INIT = 16'h0a88;
    SB_LUT4 led_counter_1186_1260_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_68), .I3(n10177), .O(n124)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4460_3_lut (.I0(\REG.mem_55_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n10), .I3(GND_net), .O(n5843));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4461_3_lut (.I0(\REG.mem_55_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n10), .I3(GND_net), .O(n5844));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4462_3_lut (.I0(\REG.mem_55_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n10), .I3(GND_net), .O(n5845));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4463_3_lut (.I0(\REG.mem_55_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n10), .I3(GND_net), .O(n5846));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4464_3_lut (.I0(\REG.mem_55_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n10), .I3(GND_net), .O(n5847));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4465_3_lut (.I0(\REG.mem_55_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n10), .I3(GND_net), .O(n5848));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4466_3_lut (.I0(\REG.mem_55_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n10), .I3(GND_net), .O(n5849));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4466_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4467_3_lut (.I0(\REG.mem_55_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n10), .I3(GND_net), .O(n5850));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4468_3_lut (.I0(\REG.mem_55_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n10), .I3(GND_net), .O(n5851));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4469_3_lut (.I0(\REG.mem_55_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n10), .I3(GND_net), .O(n5852));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6023_1_lut (.I0(n1774), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n7386));   // src/timing_controller.v(51[11:16])
    defparam i6023_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4470_3_lut (.I0(\REG.mem_55_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n10), .I3(GND_net), .O(n5853));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4471_3_lut (.I0(\REG.mem_55_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n10), .I3(GND_net), .O(n5854));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4472_3_lut (.I0(\REG.mem_55_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n10), .I3(GND_net), .O(n5855));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4473_3_lut (.I0(\REG.mem_55_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n10), .I3(GND_net), .O(n5856));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4474_3_lut (.I0(\REG.mem_55_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n10), .I3(GND_net), .O(n5857));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4475_3_lut (.I0(\REG.mem_55_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n10), .I3(GND_net), .O(n5858));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4476_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[6]), .I2(GND_net), 
            .I3(GND_net), .O(n5859));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4476_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4477_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5860));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4477_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4478_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5861));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4478_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4479_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5862));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4479_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4480_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5863));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4480_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4481_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5864));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4481_2_lut.LUT_INIT = 16'h4444;
    SB_DFF even_byte_flag_89 (.Q(even_byte_flag), .C(SLM_CLK_c), .D(n2944));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 i4502_3_lut (.I0(\REG.mem_57_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n8_adj_59), .I3(GND_net), .O(n5885));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4504_3_lut (.I0(\REG.mem_57_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n8_adj_59), .I3(GND_net), .O(n5887));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4505_3_lut (.I0(\REG.mem_57_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n8_adj_59), .I3(GND_net), .O(n5888));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4506_3_lut (.I0(\REG.mem_57_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n8_adj_59), .I3(GND_net), .O(n5889));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4507_3_lut (.I0(\REG.mem_57_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n8_adj_59), .I3(GND_net), .O(n5890));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4508_3_lut (.I0(\REG.mem_57_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n8_adj_59), .I3(GND_net), .O(n5891));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4509_3_lut (.I0(\REG.mem_57_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n8_adj_59), .I3(GND_net), .O(n5892));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4509_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4510_3_lut (.I0(\REG.mem_57_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n8_adj_59), .I3(GND_net), .O(n5893));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4511_3_lut (.I0(\REG.mem_57_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n8_adj_59), .I3(GND_net), .O(n5894));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4512_3_lut (.I0(\REG.mem_57_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n8_adj_59), .I3(GND_net), .O(n5895));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4513_3_lut (.I0(\REG.mem_57_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n8_adj_59), .I3(GND_net), .O(n5896));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4514_3_lut (.I0(\REG.mem_57_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n8_adj_59), .I3(GND_net), .O(n5897));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4515_3_lut (.I0(\REG.mem_57_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n8_adj_59), .I3(GND_net), .O(n5898));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4516_3_lut (.I0(\REG.mem_57_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n8_adj_59), .I3(GND_net), .O(n5899));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4517_3_lut (.I0(\REG.mem_57_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n8_adj_59), .I3(GND_net), .O(n5900));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4518_3_lut (.I0(\REG.mem_57_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n8_adj_59), .I3(GND_net), .O(n5901));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3931_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[5]), .I2(\mem_LUT.data_raw_r [5]), 
            .I3(n4459), .O(n5314));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i3931_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i3928_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[4]), .I2(\mem_LUT.data_raw_r [4]), 
            .I3(n4459), .O(n5311));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i3928_4_lut.LUT_INIT = 16'h5044;
    SB_DFF tx_data_byte_r_i0_i1 (.Q(tx_data_byte[1]), .C(SLM_CLK_c), .D(n4860));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_data_byte_r_i0_i2 (.Q(tx_data_byte[2]), .C(SLM_CLK_c), .D(n4859));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_data_byte_r_i0_i3 (.Q(tx_data_byte[3]), .C(SLM_CLK_c), .D(n4855));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_data_byte_r_i0_i4 (.Q(tx_data_byte[4]), .C(SLM_CLK_c), .D(n4845));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 i4538_2_lut (.I0(reset_per_frame), .I1(rd_addr_nxt_c_6__N_498[5]), 
            .I2(GND_net), .I3(GND_net), .O(n5921));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i4538_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4540_2_lut (.I0(reset_per_frame), .I1(rd_addr_nxt_c_6__N_498[3]), 
            .I2(GND_net), .I3(GND_net), .O(n5923));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i4540_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4541_2_lut (.I0(reset_per_frame), .I1(rd_addr_nxt_c_6__N_498[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5924));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i4541_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4543_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[6]), .I2(GND_net), 
            .I3(GND_net), .O(n5926));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4543_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4544_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5927));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4544_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4545_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5928));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4545_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4562_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5945));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4562_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4563_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5946));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4563_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4564_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5947));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4564_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4565_2_lut (.I0(reset_per_frame), .I1(rd_addr_r[6]), .I2(GND_net), 
            .I3(GND_net), .O(n5948));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4565_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4566_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5949));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4566_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4567_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5950));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4567_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4568_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5951));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4568_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4569_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5952));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4569_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4570_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5953));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4570_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4587_3_lut (.I0(tx_data_byte[5]), .I1(pc_data_rx[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5970));   // src/top.v(1074[8] 1141[4])
    defparam i4587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4485_4_lut_4_lut_4_lut (.I0(wr_fifo_en_w), .I1(reset_all_w), 
            .I2(wr_addr_r_adj_118[0]), .I3(wr_addr_r_adj_118[1]), .O(n5868));
    defparam i4485_4_lut_4_lut_4_lut.LUT_INIT = 16'h1320;
    SB_LUT4 i4606_4_lut_4_lut (.I0(wr_fifo_en_w), .I1(reset_all_w), .I2(wr_addr_p1_w_adj_120[2]), 
            .I3(wr_addr_r_adj_118[2]), .O(n5989));
    defparam i4606_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_DFFSR multi_byte_spi_trans_flag_r_86 (.Q(multi_byte_spi_trans_flag_r), 
            .C(SLM_CLK_c), .D(multi_byte_spi_trans_flag_r_N_72), .R(n4661));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 i3_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[3]), 
            .I3(n10871), .O(n10808));   // src/timing_controller.v(62[5] 131[12])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i10313_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(n10831), .O(n12063));   // src/timing_controller.v(62[5] 131[12])
    defparam i10313_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i6227_2_lut_3_lut (.I0(state[1]), .I1(state[0]), .I2(n63), 
            .I3(GND_net), .O(n7590));   // src/timing_controller.v(62[5] 131[12])
    defparam i6227_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i3_4_lut (.I0(reset_clk_counter[0]), .I1(reset_clk_counter[2]), 
            .I2(reset_clk_counter[3]), .I3(reset_clk_counter[1]), .O(reset_all_w_N_61));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF tx_data_byte_r_i0_i0 (.Q(tx_data_byte[0]), .C(SLM_CLK_c), .D(n4824));   // src/top.v(1074[8] 1141[4])
    SB_CARRY led_counter_1186_1260_add_4_8 (.CI(n10177), .I0(GND_net), .I1(n19_adj_68), 
            .CO(n10178));
    SB_DFF fifo_read_cmd_80 (.Q(fifo_read_cmd), .C(SLM_CLK_c), .D(start_tx_N_64));   // src/top.v(910[8] 928[4])
    SB_LUT4 led_counter_1186_1260_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_67), .I3(n10176), .O(n125)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_7 (.CI(n10176), .I0(GND_net), .I1(n20_adj_67), 
            .CO(n10177));
    SB_LUT4 led_counter_1186_1260_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_66), .I3(n10175), .O(n126)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3507_3_lut (.I0(r_Tx_Data[0]), .I1(fifo_temp_output[0]), .I2(n3794), 
            .I3(GND_net), .O(n4890));   // src/uart_tx.v(38[10] 141[8])
    defparam i3507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3505_3_lut (.I0(rx_shift_reg[1]), .I1(rx_shift_reg[0]), .I2(n4312), 
            .I3(GND_net), .O(n4888));   // src/spi.v(76[8] 221[4])
    defparam i3505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4058_3_lut (.I0(\REG.mem_31_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n34), .I3(GND_net), .O(n5441));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4057_3_lut (.I0(\REG.mem_31_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n34), .I3(GND_net), .O(n5440));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4056_3_lut (.I0(\REG.mem_31_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n34), .I3(GND_net), .O(n5439));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4055_3_lut (.I0(\REG.mem_31_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n34), .I3(GND_net), .O(n5438));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4054_3_lut (.I0(\REG.mem_31_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n34), .I3(GND_net), .O(n5437));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4053_3_lut (.I0(\REG.mem_31_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n34), .I3(GND_net), .O(n5436));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4052_3_lut (.I0(\REG.mem_31_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n34), .I3(GND_net), .O(n5435));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4051_3_lut (.I0(\REG.mem_31_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n34), .I3(GND_net), .O(n5434));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4050_3_lut (.I0(\REG.mem_31_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n34), .I3(GND_net), .O(n5433));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4049_3_lut (.I0(\REG.mem_31_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n34), .I3(GND_net), .O(n5432));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4048_3_lut (.I0(\REG.mem_31_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n34), .I3(GND_net), .O(n5431));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4047_3_lut (.I0(\REG.mem_31_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n34), .I3(GND_net), .O(n5430));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4046_3_lut (.I0(\REG.mem_31_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n34), .I3(GND_net), .O(n5429));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4045_3_lut (.I0(\REG.mem_31_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n34), .I3(GND_net), .O(n5428));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4044_3_lut (.I0(\REG.mem_31_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n34), .I3(GND_net), .O(n5427));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4043_3_lut (.I0(\REG.mem_31_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n34), .I3(GND_net), .O(n5426));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_76));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3500_3_lut (.I0(rx_shift_reg[2]), .I1(rx_shift_reg[1]), .I2(n4312), 
            .I3(GND_net), .O(n4883));   // src/spi.v(76[8] 221[4])
    defparam i3500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3962_3_lut (.I0(\REG.mem_25_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n40), .I3(GND_net), .O(n5345));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3961_3_lut (.I0(\REG.mem_25_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n40), .I3(GND_net), .O(n5344));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3960_3_lut (.I0(\REG.mem_25_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n40), .I3(GND_net), .O(n5343));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3959_3_lut (.I0(\REG.mem_25_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n40), .I3(GND_net), .O(n5342));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3958_3_lut (.I0(\REG.mem_25_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n40), .I3(GND_net), .O(n5341));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3957_3_lut (.I0(\REG.mem_25_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n40), .I3(GND_net), .O(n5340));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3956_3_lut (.I0(\REG.mem_25_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n40), .I3(GND_net), .O(n5339));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3955_3_lut (.I0(\REG.mem_25_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n40), .I3(GND_net), .O(n5338));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3954_3_lut (.I0(\REG.mem_25_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n40), .I3(GND_net), .O(n5337));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3953_3_lut (.I0(\REG.mem_25_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n40), .I3(GND_net), .O(n5336));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3952_3_lut (.I0(\REG.mem_25_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n40), .I3(GND_net), .O(n5335));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3951_3_lut (.I0(\REG.mem_25_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n40), .I3(GND_net), .O(n5334));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3950_3_lut (.I0(\REG.mem_25_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n40), .I3(GND_net), .O(n5333));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3949_3_lut (.I0(\REG.mem_25_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n40), .I3(GND_net), .O(n5332));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3948_3_lut (.I0(\REG.mem_25_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n40), .I3(GND_net), .O(n5331));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3947_3_lut (.I0(\REG.mem_25_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n40), .I3(GND_net), .O(n5330));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3923_3_lut (.I0(\REG.mem_23_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n42), .I3(GND_net), .O(n5306));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3922_3_lut (.I0(\REG.mem_23_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n42), .I3(GND_net), .O(n5305));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3921_3_lut (.I0(\REG.mem_23_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n42), .I3(GND_net), .O(n5304));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3920_3_lut (.I0(\REG.mem_23_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n42), .I3(GND_net), .O(n5303));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3919_3_lut (.I0(\REG.mem_23_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n42), .I3(GND_net), .O(n5302));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3918_3_lut (.I0(\REG.mem_23_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n42), .I3(GND_net), .O(n5301));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3917_3_lut (.I0(\REG.mem_23_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n42), .I3(GND_net), .O(n5300));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3916_3_lut (.I0(\REG.mem_23_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n42), .I3(GND_net), .O(n5299));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3915_3_lut (.I0(\REG.mem_23_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n42), .I3(GND_net), .O(n5298));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3914_3_lut (.I0(\REG.mem_23_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n42), .I3(GND_net), .O(n5297));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3913_3_lut (.I0(\REG.mem_23_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n42), .I3(GND_net), .O(n5296));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3912_3_lut (.I0(\REG.mem_23_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n42), .I3(GND_net), .O(n5295));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3911_3_lut (.I0(\REG.mem_23_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n42), .I3(GND_net), .O(n5294));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3910_3_lut (.I0(\REG.mem_23_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n42), .I3(GND_net), .O(n5293));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3909_3_lut (.I0(\REG.mem_23_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n42), .I3(GND_net), .O(n5292));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3907_3_lut (.I0(\REG.mem_23_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n42), .I3(GND_net), .O(n5290));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3841_3_lut (.I0(\REG.mem_18_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n47), .I3(GND_net), .O(n5224));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3840_3_lut (.I0(\REG.mem_18_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n47), .I3(GND_net), .O(n5223));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3839_3_lut (.I0(\REG.mem_18_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n47), .I3(GND_net), .O(n5222));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3838_3_lut (.I0(\REG.mem_18_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n47), .I3(GND_net), .O(n5221));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3837_3_lut (.I0(\REG.mem_18_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n47), .I3(GND_net), .O(n5220));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3836_3_lut (.I0(\REG.mem_18_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n47), .I3(GND_net), .O(n5219));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3835_3_lut (.I0(\REG.mem_18_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n47), .I3(GND_net), .O(n5218));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3834_3_lut (.I0(\REG.mem_18_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n47), .I3(GND_net), .O(n5217));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3833_3_lut (.I0(\REG.mem_18_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n47), .I3(GND_net), .O(n5216));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3832_3_lut (.I0(\REG.mem_18_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n47), .I3(GND_net), .O(n5215));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3831_3_lut (.I0(\REG.mem_18_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n47), .I3(GND_net), .O(n5214));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3830_3_lut (.I0(\REG.mem_18_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n47), .I3(GND_net), .O(n5213));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3829_3_lut (.I0(\REG.mem_18_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n47), .I3(GND_net), .O(n5212));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3828_3_lut (.I0(\REG.mem_18_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n47), .I3(GND_net), .O(n5211));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3827_3_lut (.I0(\REG.mem_18_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n47), .I3(GND_net), .O(n5210));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3826_3_lut (.I0(\REG.mem_18_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n47), .I3(GND_net), .O(n5209));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3278_1_lut_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n4661));   // src/top.v(1074[8] 1141[4])
    defparam i3278_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(rd_fifo_en_prev_r), .I1(fifo_read_cmd), 
            .I2(is_fifo_empty_flag), .I3(reset_all_w), .O(n4459));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hffae;
    SB_LUT4 i3495_2_lut_3_lut (.I0(reset_all_w), .I1(fifo_read_cmd), .I2(is_fifo_empty_flag), 
            .I3(GND_net), .O(n4878));   // src/fifo_quad_word_mod.v(353[29] 363[32])
    defparam i3495_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1590_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n2944));   // src/top.v(1074[8] 1141[4])
    defparam i1590_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3506_4_lut_4_lut (.I0(tx_uart_active_flag), .I1(r_SM_Main_adj_95[1]), 
            .I2(r_SM_Main_adj_95[2]), .I3(n10805), .O(n4889));   // src/uart_tx.v(38[10] 141[8])
    defparam i3506_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i3809_3_lut (.I0(r_Tx_Data[1]), .I1(fifo_temp_output[1]), .I2(n3794), 
            .I3(GND_net), .O(n5192));   // src/uart_tx.v(38[10] 141[8])
    defparam i3809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3808_3_lut (.I0(r_Tx_Data[2]), .I1(fifo_temp_output[2]), .I2(n3794), 
            .I3(GND_net), .O(n5191));   // src/uart_tx.v(38[10] 141[8])
    defparam i3808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3807_3_lut (.I0(r_Tx_Data[3]), .I1(fifo_temp_output[3]), .I2(n3794), 
            .I3(GND_net), .O(n5190));   // src/uart_tx.v(38[10] 141[8])
    defparam i3807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3806_3_lut (.I0(r_Tx_Data[4]), .I1(fifo_temp_output[4]), .I2(n3794), 
            .I3(GND_net), .O(n5189));   // src/uart_tx.v(38[10] 141[8])
    defparam i3806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3805_3_lut (.I0(\REG.mem_16_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n49), .I3(GND_net), .O(n5188));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3804_3_lut (.I0(r_Tx_Data[5]), .I1(fifo_temp_output[5]), .I2(n3794), 
            .I3(GND_net), .O(n5187));   // src/uart_tx.v(38[10] 141[8])
    defparam i3804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3803_3_lut (.I0(\REG.mem_16_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n49), .I3(GND_net), .O(n5186));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3802_3_lut (.I0(\REG.mem_16_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n49), .I3(GND_net), .O(n5185));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3801_3_lut (.I0(\REG.mem_16_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n49), .I3(GND_net), .O(n5184));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3800_3_lut (.I0(\REG.mem_16_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n49), .I3(GND_net), .O(n5183));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3799_3_lut (.I0(\REG.mem_16_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n49), .I3(GND_net), .O(n5182));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3798_3_lut (.I0(\REG.mem_16_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n49), .I3(GND_net), .O(n5181));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3797_3_lut (.I0(\REG.mem_16_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n49), .I3(GND_net), .O(n5180));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3796_3_lut (.I0(\REG.mem_16_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n49), .I3(GND_net), .O(n5179));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3795_3_lut (.I0(\REG.mem_16_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n49), .I3(GND_net), .O(n5178));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3794_3_lut (.I0(\REG.mem_16_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n49), .I3(GND_net), .O(n5177));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3793_3_lut (.I0(\REG.mem_16_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n49), .I3(GND_net), .O(n5176));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1601_2_lut_3_lut_4_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(reset_all_w), .I3(wr_addr_r_adj_118[0]), .O(n8));
    defparam i1601_2_lut_3_lut_4_lut.LUT_INIT = 16'h0df2;
    SB_LUT4 i3792_3_lut (.I0(\REG.mem_16_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n49), .I3(GND_net), .O(n5175));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3791_3_lut (.I0(\REG.mem_16_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n49), .I3(GND_net), .O(n5174));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3790_3_lut (.I0(\REG.mem_16_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n49), .I3(GND_net), .O(n5173));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3789_3_lut (.I0(\REG.mem_16_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n49), .I3(GND_net), .O(n5172));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3788_3_lut (.I0(r_Tx_Data[6]), .I1(fifo_temp_output[6]), .I2(n3794), 
            .I3(GND_net), .O(n5171));   // src/uart_tx.v(38[10] 141[8])
    defparam i3788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3787_3_lut (.I0(r_Tx_Data[7]), .I1(fifo_temp_output[7]), .I2(n3794), 
            .I3(GND_net), .O(n5170));   // src/uart_tx.v(38[10] 141[8])
    defparam i3787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3786_3_lut (.I0(\REG.mem_15_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n50), .I3(GND_net), .O(n5169));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3785_3_lut (.I0(\REG.mem_15_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n50), .I3(GND_net), .O(n5168));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3784_3_lut (.I0(\REG.mem_15_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n50), .I3(GND_net), .O(n5167));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3783_3_lut (.I0(\REG.mem_15_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n50), .I3(GND_net), .O(n5166));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3782_3_lut (.I0(\REG.mem_15_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n50), .I3(GND_net), .O(n5165));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3781_3_lut (.I0(\REG.mem_15_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n50), .I3(GND_net), .O(n5164));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3780_3_lut (.I0(\REG.mem_15_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n50), .I3(GND_net), .O(n5163));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3779_3_lut (.I0(\REG.mem_15_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n50), .I3(GND_net), .O(n5162));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3778_3_lut (.I0(\REG.mem_15_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n50), .I3(GND_net), .O(n5161));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3777_3_lut (.I0(\REG.mem_15_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n50), .I3(GND_net), .O(n5160));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3776_3_lut (.I0(\REG.mem_15_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n50), .I3(GND_net), .O(n5159));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3775_3_lut (.I0(\REG.mem_15_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n50), .I3(GND_net), .O(n5158));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3774_3_lut (.I0(\REG.mem_15_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n50), .I3(GND_net), .O(n5157));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3773_3_lut (.I0(\REG.mem_15_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n50), .I3(GND_net), .O(n5156));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3772_3_lut (.I0(\REG.mem_15_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n50), .I3(GND_net), .O(n5155));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3771_3_lut (.I0(\REG.mem_15_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n50), .I3(GND_net), .O(n5154));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3770_3_lut (.I0(\REG.mem_14_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n51), .I3(GND_net), .O(n5153));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3770_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3769_3_lut (.I0(\REG.mem_14_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n51), .I3(GND_net), .O(n5152));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3768_3_lut (.I0(\REG.mem_14_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n51), .I3(GND_net), .O(n5151));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3767_3_lut (.I0(\REG.mem_14_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n51), .I3(GND_net), .O(n5150));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3766_3_lut (.I0(\REG.mem_14_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n51), .I3(GND_net), .O(n5149));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3765_3_lut (.I0(\REG.mem_14_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n51), .I3(GND_net), .O(n5148));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3764_3_lut (.I0(\REG.mem_14_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n51), .I3(GND_net), .O(n5147));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3763_3_lut (.I0(\REG.mem_14_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n51), .I3(GND_net), .O(n5146));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3762_3_lut (.I0(\REG.mem_14_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n51), .I3(GND_net), .O(n5145));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3761_3_lut (.I0(\REG.mem_14_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n51), .I3(GND_net), .O(n5144));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3760_3_lut (.I0(\REG.mem_14_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n51), .I3(GND_net), .O(n5143));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3759_3_lut (.I0(\REG.mem_14_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n51), .I3(GND_net), .O(n5142));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3758_3_lut (.I0(\REG.mem_14_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n51), .I3(GND_net), .O(n5141));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3757_3_lut (.I0(\REG.mem_14_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n51), .I3(GND_net), .O(n5140));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3756_3_lut (.I0(\REG.mem_14_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n51), .I3(GND_net), .O(n5139));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3755_3_lut (.I0(\REG.mem_14_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n51), .I3(GND_net), .O(n5138));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3754_3_lut (.I0(\REG.mem_13_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n52), .I3(GND_net), .O(n5137));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3753_3_lut (.I0(\REG.mem_13_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n52), .I3(GND_net), .O(n5136));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3752_3_lut (.I0(\REG.mem_13_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n52), .I3(GND_net), .O(n5135));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3751_3_lut (.I0(\REG.mem_13_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n52), .I3(GND_net), .O(n5134));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3750_3_lut (.I0(\REG.mem_13_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n52), .I3(GND_net), .O(n5133));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3494_3_lut (.I0(rx_shift_reg[3]), .I1(rx_shift_reg[2]), .I2(n4312), 
            .I3(GND_net), .O(n4877));   // src/spi.v(76[8] 221[4])
    defparam i3494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3749_3_lut (.I0(\REG.mem_13_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n52), .I3(GND_net), .O(n5132));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3748_3_lut (.I0(\REG.mem_13_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n52), .I3(GND_net), .O(n5131));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3747_3_lut (.I0(\REG.mem_13_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n52), .I3(GND_net), .O(n5130));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3746_3_lut (.I0(\REG.mem_13_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n52), .I3(GND_net), .O(n5129));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3745_3_lut (.I0(\REG.mem_13_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n52), .I3(GND_net), .O(n5128));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3744_3_lut (.I0(\REG.mem_13_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n52), .I3(GND_net), .O(n5127));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3743_3_lut (.I0(\REG.mem_13_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n52), .I3(GND_net), .O(n5126));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3742_3_lut (.I0(\REG.mem_13_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n52), .I3(GND_net), .O(n5125));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3741_3_lut (.I0(\REG.mem_13_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n52), .I3(GND_net), .O(n5124));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3740_3_lut (.I0(\REG.mem_13_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n52), .I3(GND_net), .O(n5123));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3739_3_lut (.I0(\REG.mem_13_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n52), .I3(GND_net), .O(n5122));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3738_3_lut (.I0(\REG.mem_12_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n53), .I3(GND_net), .O(n5121));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3737_3_lut (.I0(\REG.mem_12_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n53), .I3(GND_net), .O(n5120));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3736_3_lut (.I0(\REG.mem_12_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n53), .I3(GND_net), .O(n5119));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3735_3_lut (.I0(\REG.mem_12_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n53), .I3(GND_net), .O(n5118));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3734_3_lut (.I0(\REG.mem_12_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n53), .I3(GND_net), .O(n5117));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3733_3_lut (.I0(\REG.mem_12_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n53), .I3(GND_net), .O(n5116));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3486_3_lut (.I0(rx_shift_reg[4]), .I1(rx_shift_reg[3]), .I2(n4312), 
            .I3(GND_net), .O(n4869));   // src/spi.v(76[8] 221[4])
    defparam i3486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3732_3_lut (.I0(\REG.mem_12_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n53), .I3(GND_net), .O(n5115));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3731_3_lut (.I0(\REG.mem_12_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n53), .I3(GND_net), .O(n5114));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3730_3_lut (.I0(\REG.mem_12_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n53), .I3(GND_net), .O(n5113));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3729_3_lut (.I0(\REG.mem_12_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n53), .I3(GND_net), .O(n5112));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3728_3_lut (.I0(\REG.mem_12_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n53), .I3(GND_net), .O(n5111));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3727_3_lut (.I0(\REG.mem_12_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n53), .I3(GND_net), .O(n5110));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3726_3_lut (.I0(\REG.mem_12_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n53), .I3(GND_net), .O(n5109));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3725_3_lut (.I0(\REG.mem_12_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n53), .I3(GND_net), .O(n5108));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3724_3_lut (.I0(\REG.mem_12_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n53), .I3(GND_net), .O(n5107));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3724_3_lut.LUT_INIT = 16'hcaca;
    fifo_dc_32_lut_gen2 fifo_dc_32_lut_gen_inst (.\rd_addr_r[0] (rd_addr_r[0]), 
            .\REG.mem_14_5 (\REG.mem_14_5 ), .\REG.mem_15_5 (\REG.mem_15_5 ), 
            .\dc32_fifo_data_in[6] (dc32_fifo_data_in[6]), .dc32_fifo_almost_full(dc32_fifo_almost_full), 
            .FIFO_CLK_c(FIFO_CLK_c), .reset_per_frame(reset_per_frame), 
            .\REG.mem_13_5 (\REG.mem_13_5 ), .\REG.mem_12_5 (\REG.mem_12_5 ), 
            .\dc32_fifo_data_in[5] (dc32_fifo_data_in[5]), .\dc32_fifo_data_in[4] (dc32_fifo_data_in[4]), 
            .\REG.mem_31_0 (\REG.mem_31_0 ), .GND_net(GND_net), .\dc32_fifo_data_in[3] (dc32_fifo_data_in[3]), 
            .\REG.mem_55_13 (\REG.mem_55_13 ), .\dc32_fifo_data_in[2] (dc32_fifo_data_in[2]), 
            .\REG.mem_38_7 (\REG.mem_38_7 ), .\REG.mem_39_7 (\REG.mem_39_7 ), 
            .\REG.mem_36_7 (\REG.mem_36_7 ), .\REG.mem_37_7 (\REG.mem_37_7 ), 
            .\REG.mem_16_8 (\REG.mem_16_8 ), .\REG.mem_18_8 (\REG.mem_18_8 ), 
            .\REG.mem_3_13 (\REG.mem_3_13 ), .\REG.mem_57_6 (\REG.mem_57_6 ), 
            .\dc32_fifo_data_in[1] (dc32_fifo_data_in[1]), .\REG.mem_63_11 (\REG.mem_63_11 ), 
            .\dc32_fifo_data_in[0] (dc32_fifo_data_in[0]), .\REG.mem_35_0 (\REG.mem_35_0 ), 
            .t_rd_fifo_en_w(t_rd_fifo_en_w), .\REG.out_raw[0] (\REG.out_raw [0]), 
            .SLM_CLK_c(SLM_CLK_c), .\REG.mem_55_10 (\REG.mem_55_10 ), .n62(n62), 
            .n30(n30), .\REG.mem_31_3 (\REG.mem_31_3 ), .\REG.mem_48_7 (\REG.mem_48_7 ), 
            .\REG.mem_50_7 (\REG.mem_50_7 ), .\REG.mem_55_7 (\REG.mem_55_7 ), 
            .\REG.mem_48_10 (\REG.mem_48_10 ), .\REG.mem_50_10 (\REG.mem_50_10 ), 
            .wr_grey_sync_r({wr_grey_sync_r}), .\wr_addr_nxt_c[5] (wr_addr_nxt_c[5]), 
            .\REG.mem_23_8 (\REG.mem_23_8 ), .\REG.mem_25_5 (\REG.mem_25_5 ), 
            .\rd_grey_sync_r[0] (rd_grey_sync_r[0]), .\REG.mem_25_15 (\REG.mem_25_15 ), 
            .\REG.mem_14_12 (\REG.mem_14_12 ), .\REG.mem_15_12 (\REG.mem_15_12 ), 
            .DEBUG_3_c(DEBUG_3_c), .\REG.mem_13_12 (\REG.mem_13_12 ), .\REG.mem_12_12 (\REG.mem_12_12 ), 
            .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .dc32_fifo_almost_empty(dc32_fifo_almost_empty), .\REG.mem_6_1 (\REG.mem_6_1 ), 
            .\REG.mem_7_1 (\REG.mem_7_1 ), .\REG.mem_5_1 (\REG.mem_5_1 ), 
            .\REG.mem_4_1 (\REG.mem_4_1 ), .\REG.mem_57_9 (\REG.mem_57_9 ), 
            .\REG.mem_35_3 (\REG.mem_35_3 ), .\REG.mem_46_1 (\REG.mem_46_1 ), 
            .\REG.mem_47_1 (\REG.mem_47_1 ), .\REG.mem_45_1 (\REG.mem_45_1 ), 
            .\REG.mem_44_1 (\REG.mem_44_1 ), .\REG.mem_25_2 (\REG.mem_25_2 ), 
            .\dc32_fifo_data_in[15] (dc32_fifo_data_in[15]), .\dc32_fifo_data_in[14] (dc32_fifo_data_in[14]), 
            .\dc32_fifo_data_in[13] (dc32_fifo_data_in[13]), .\REG.mem_3_11 (\REG.mem_3_11 ), 
            .\REG.mem_31_2 (\REG.mem_31_2 ), .\REG.mem_50_12 (\REG.mem_50_12 ), 
            .\dc32_fifo_data_in[12] (dc32_fifo_data_in[12]), .\REG.mem_6_11 (\REG.mem_6_11 ), 
            .\REG.mem_7_11 (\REG.mem_7_11 ), .\REG.mem_5_11 (\REG.mem_5_11 ), 
            .\REG.mem_4_11 (\REG.mem_4_11 ), .\dc32_fifo_data_in[11] (dc32_fifo_data_in[11]), 
            .\REG.mem_48_12 (\REG.mem_48_12 ), .\REG.mem_3_4 (\REG.mem_3_4 ), 
            .\REG.mem_14_8 (\REG.mem_14_8 ), .\REG.mem_15_8 (\REG.mem_15_8 ), 
            .\REG.mem_8_14 (\REG.mem_8_14 ), .\REG.mem_9_14 (\REG.mem_9_14 ), 
            .\dc32_fifo_data_in[10] (dc32_fifo_data_in[10]), .\REG.mem_10_14 (\REG.mem_10_14 ), 
            .\REG.mem_11_14 (\REG.mem_11_14 ), .\REG.mem_63_6 (\REG.mem_63_6 ), 
            .\REG.mem_13_8 (\REG.mem_13_8 ), .\REG.mem_12_8 (\REG.mem_12_8 ), 
            .\REG.mem_14_14 (\REG.mem_14_14 ), .\REG.mem_15_14 (\REG.mem_15_14 ), 
            .\dc32_fifo_data_in[9] (dc32_fifo_data_in[9]), .\dc32_fifo_data_in[8] (dc32_fifo_data_in[8]), 
            .\REG.mem_3_1 (\REG.mem_3_1 ), .\dc32_fifo_data_in[7] (dc32_fifo_data_in[7]), 
            .\REG.mem_12_14 (\REG.mem_12_14 ), .\REG.mem_13_14 (\REG.mem_13_14 ), 
            .\REG.mem_42_8 (\REG.mem_42_8 ), .\REG.mem_43_8 (\REG.mem_43_8 ), 
            .\REG.mem_41_8 (\REG.mem_41_8 ), .\REG.mem_40_8 (\REG.mem_40_8 ), 
            .\REG.mem_18_12 (\REG.mem_18_12 ), .\REG.mem_16_12 (\REG.mem_16_12 ), 
            .\REG.mem_31_15 (\REG.mem_31_15 ), .\REG.mem_38_3 (\REG.mem_38_3 ), 
            .\REG.mem_39_3 (\REG.mem_39_3 ), .\REG.mem_37_3 (\REG.mem_37_3 ), 
            .\REG.mem_36_3 (\REG.mem_36_3 ), .\REG.mem_42_3 (\REG.mem_42_3 ), 
            .\REG.mem_43_3 (\REG.mem_43_3 ), .\REG.mem_14_7 (\REG.mem_14_7 ), 
            .\REG.mem_15_7 (\REG.mem_15_7 ), .\REG.mem_13_7 (\REG.mem_13_7 ), 
            .\REG.mem_12_7 (\REG.mem_12_7 ), .\REG.mem_41_3 (\REG.mem_41_3 ), 
            .\REG.mem_40_3 (\REG.mem_40_3 ), .\REG.mem_57_0 (\REG.mem_57_0 ), 
            .\REG.mem_10_11 (\REG.mem_10_11 ), .\REG.mem_11_11 (\REG.mem_11_11 ), 
            .\REG.mem_9_11 (\REG.mem_9_11 ), .\REG.mem_8_11 (\REG.mem_8_11 ), 
            .\REG.mem_63_12 (\REG.mem_63_12 ), .\REG.mem_55_12 (\REG.mem_55_12 ), 
            .\REG.mem_35_15 (\REG.mem_35_15 ), .\REG.mem_3_15 (\REG.mem_3_15 ), 
            .\wr_addr_nxt_c[3] (wr_addr_nxt_c[3]), .\REG.mem_50_9 (\REG.mem_50_9 ), 
            .\REG.mem_48_9 (\REG.mem_48_9 ), .\REG.mem_46_8 (\REG.mem_46_8 ), 
            .\REG.mem_47_8 (\REG.mem_47_8 ), .\REG.mem_46_3 (\REG.mem_46_3 ), 
            .\REG.mem_47_3 (\REG.mem_47_3 ), .\REG.mem_45_8 (\REG.mem_45_8 ), 
            .\REG.mem_44_8 (\REG.mem_44_8 ), .\REG.mem_16_2 (\REG.mem_16_2 ), 
            .\REG.mem_10_9 (\REG.mem_10_9 ), .\REG.mem_11_9 (\REG.mem_11_9 ), 
            .\REG.mem_45_3 (\REG.mem_45_3 ), .\REG.mem_44_3 (\REG.mem_44_3 ), 
            .\REG.mem_25_7 (\REG.mem_25_7 ), .\REG.mem_23_12 (\REG.mem_23_12 ), 
            .\REG.mem_18_2 (\REG.mem_18_2 ), .\REG.mem_38_0 (\REG.mem_38_0 ), 
            .\REG.mem_39_0 (\REG.mem_39_0 ), .\REG.mem_31_13 (\REG.mem_31_13 ), 
            .\REG.mem_37_0 (\REG.mem_37_0 ), .\REG.mem_36_0 (\REG.mem_36_0 ), 
            .\REG.mem_18_6 (\REG.mem_18_6 ), .\REG.mem_16_6 (\REG.mem_16_6 ), 
            .\REG.mem_9_9 (\REG.mem_9_9 ), .\REG.mem_8_9 (\REG.mem_8_9 ), 
            .\REG.mem_50_3 (\REG.mem_50_3 ), .\REG.mem_48_3 (\REG.mem_48_3 ), 
            .\REG.mem_42_0 (\REG.mem_42_0 ), .\REG.mem_43_0 (\REG.mem_43_0 ), 
            .\REG.mem_41_0 (\REG.mem_41_0 ), .\REG.mem_40_0 (\REG.mem_40_0 ), 
            .\REG.mem_14_11 (\REG.mem_14_11 ), .\REG.mem_15_11 (\REG.mem_15_11 ), 
            .\REG.mem_13_11 (\REG.mem_13_11 ), .\REG.mem_12_11 (\REG.mem_12_11 ), 
            .\REG.mem_38_5 (\REG.mem_38_5 ), .\REG.mem_39_5 (\REG.mem_39_5 ), 
            .\REG.mem_37_5 (\REG.mem_37_5 ), .\REG.mem_36_5 (\REG.mem_36_5 ), 
            .\REG.mem_57_13 (\REG.mem_57_13 ), .n6121(n6121), .VCC_net(VCC_net), 
            .\fifo_data_out[2] (fifo_data_out[2]), .n6118(n6118), .\fifo_data_out[1] (fifo_data_out[1]), 
            .\REG.mem_50_1 (\REG.mem_50_1 ), .\REG.mem_6_9 (\REG.mem_6_9 ), 
            .\REG.mem_7_9 (\REG.mem_7_9 ), .\REG.mem_48_1 (\REG.mem_48_1 ), 
            .n10556(n10556), .\fifo_data_out[3] (fifo_data_out[3]), .n10562(n10562), 
            .\fifo_data_out[4] (fifo_data_out[4]), .\REG.mem_18_11 (\REG.mem_18_11 ), 
            .\REG.mem_16_11 (\REG.mem_16_11 ), .\REG.mem_5_9 (\REG.mem_5_9 ), 
            .\REG.mem_4_9 (\REG.mem_4_9 ), .n10564(n10564), .\fifo_data_out[5] (fifo_data_out[5]), 
            .n10566(n10566), .\fifo_data_out[6] (fifo_data_out[6]), .n10568(n10568), 
            .\fifo_data_out[7] (fifo_data_out[7]), .n10570(n10570), .\fifo_data_out[8] (fifo_data_out[8]), 
            .n10572(n10572), .\fifo_data_out[9] (fifo_data_out[9]), .n10574(n10574), 
            .\fifo_data_out[10] (fifo_data_out[10]), .n10576(n10576), .\fifo_data_out[11] (fifo_data_out[11]), 
            .\REG.mem_31_5 (\REG.mem_31_5 ), .n6085(n6085), .\fifo_data_out[0] (fifo_data_out[0]), 
            .\REG.mem_25_12 (\REG.mem_25_12 ), .\REG.mem_38_13 (\REG.mem_38_13 ), 
            .\REG.mem_39_13 (\REG.mem_39_13 ), .n10578(n10578), .\fifo_data_out[12] (fifo_data_out[12]), 
            .n10580(n10580), .\fifo_data_out[13] (fifo_data_out[13]), .\rd_addr_r[6] (rd_addr_r[6]), 
            .\REG.mem_6_15 (\REG.mem_6_15 ), .\REG.mem_7_15 (\REG.mem_7_15 ), 
            .n6045(n6045), .n6043(n6043), .\REG.mem_5_15 (\REG.mem_5_15 ), 
            .\REG.mem_4_15 (\REG.mem_4_15 ), .\REG.mem_35_13 (\REG.mem_35_13 ), 
            .n6024(n6024), .n6021(n6021), .\REG.mem_63_15 (\REG.mem_63_15 ), 
            .n6020(n6020), .\REG.mem_63_14 (\REG.mem_63_14 ), .n6019(n6019), 
            .\REG.mem_63_13 (\REG.mem_63_13 ), .n6018(n6018), .n6017(n6017), 
            .n6016(n6016), .\REG.mem_63_10 (\REG.mem_63_10 ), .n6015(n6015), 
            .\REG.mem_63_9 (\REG.mem_63_9 ), .n6014(n6014), .\REG.mem_63_8 (\REG.mem_63_8 ), 
            .n6013(n6013), .\REG.mem_63_7 (\REG.mem_63_7 ), .n6012(n6012), 
            .n6011(n6011), .\REG.mem_63_5 (\REG.mem_63_5 ), .n6010(n6010), 
            .\REG.mem_63_4 (\REG.mem_63_4 ), .n6009(n6009), .\REG.mem_63_3 (\REG.mem_63_3 ), 
            .n6008(n6008), .\REG.mem_63_2 (\REG.mem_63_2 ), .n6007(n6007), 
            .\REG.mem_63_1 (\REG.mem_63_1 ), .n6006(n6006), .\REG.mem_63_0 (\REG.mem_63_0 ), 
            .\REG.mem_25_6 (\REG.mem_25_6 ), .\REG.mem_37_13 (\REG.mem_37_13 ), 
            .\REG.mem_36_13 (\REG.mem_36_13 ), .\REG.mem_57_4 (\REG.mem_57_4 ), 
            .\REG.mem_18_7 (\REG.mem_18_7 ), .\REG.mem_16_7 (\REG.mem_16_7 ), 
            .\REG.mem_38_15 (\REG.mem_38_15 ), .\REG.mem_39_15 (\REG.mem_39_15 ), 
            .\REG.mem_23_11 (\REG.mem_23_11 ), .\REG.mem_37_15 (\REG.mem_37_15 ), 
            .\REG.mem_36_15 (\REG.mem_36_15 ), .\REG.mem_25_11 (\REG.mem_25_11 ), 
            .\REG.mem_57_12 (\REG.mem_57_12 ), .\REG.mem_40_14 (\REG.mem_40_14 ), 
            .\REG.mem_41_14 (\REG.mem_41_14 ), .n5953(n5953), .rp_sync1_r({rp_sync1_r}), 
            .\REG.mem_42_14 (\REG.mem_42_14 ), .\REG.mem_43_14 (\REG.mem_43_14 ), 
            .\REG.mem_46_14 (\REG.mem_46_14 ), .\REG.mem_47_14 (\REG.mem_47_14 ), 
            .n5952(n5952), .n5951(n5951), .n5950(n5950), .n5949(n5949), 
            .n5948(n5948), .n5947(n5947), .n5946(n5946), .n5945(n5945), 
            .\REG.mem_55_9 (\REG.mem_55_9 ), .\REG.mem_44_14 (\REG.mem_44_14 ), 
            .\REG.mem_45_14 (\REG.mem_45_14 ), .\REG.mem_10_7 (\REG.mem_10_7 ), 
            .\REG.mem_11_7 (\REG.mem_11_7 ), .n5928(n5928), .n5927(n5927), 
            .n5926(n5926), .n5924(n5924), .n5923(n5923), .n5921(n5921), 
            .\REG.mem_9_7 (\REG.mem_9_7 ), .\REG.mem_8_7 (\REG.mem_8_7 ), 
            .\REG.mem_40_4 (\REG.mem_40_4 ), .\REG.mem_41_4 (\REG.mem_41_4 ), 
            .\REG.mem_42_4 (\REG.mem_42_4 ), .\REG.mem_43_4 (\REG.mem_43_4 ), 
            .\REG.mem_46_4 (\REG.mem_46_4 ), .\REG.mem_47_4 (\REG.mem_47_4 ), 
            .\REG.mem_44_4 (\REG.mem_44_4 ), .\REG.mem_45_4 (\REG.mem_45_4 ), 
            .n5901(n5901), .\REG.mem_57_15 (\REG.mem_57_15 ), .n5900(n5900), 
            .\REG.mem_57_14 (\REG.mem_57_14 ), .n5899(n5899), .n5898(n5898), 
            .n5897(n5897), .\REG.mem_57_11 (\REG.mem_57_11 ), .n5896(n5896), 
            .\REG.mem_57_10 (\REG.mem_57_10 ), .n5895(n5895), .n5894(n5894), 
            .\REG.mem_57_8 (\REG.mem_57_8 ), .n5893(n5893), .\REG.mem_57_7 (\REG.mem_57_7 ), 
            .n5892(n5892), .n5891(n5891), .\REG.mem_57_5 (\REG.mem_57_5 ), 
            .n5890(n5890), .n5889(n5889), .\REG.mem_57_3 (\REG.mem_57_3 ), 
            .n5888(n5888), .\REG.mem_57_2 (\REG.mem_57_2 ), .n5887(n5887), 
            .\REG.mem_57_1 (\REG.mem_57_1 ), .\REG.mem_18_1 (\REG.mem_18_1 ), 
            .\REG.mem_16_1 (\REG.mem_16_1 ), .n5885(n5885), .\REG.mem_35_8 (\REG.mem_35_8 ), 
            .\REG.mem_38_8 (\REG.mem_38_8 ), .\REG.mem_39_8 (\REG.mem_39_8 ), 
            .\REG.mem_36_8 (\REG.mem_36_8 ), .\REG.mem_37_8 (\REG.mem_37_8 ), 
            .n5864(n5864), .wp_sync1_r({wp_sync1_r}), .n5863(n5863), .n5862(n5862), 
            .n5861(n5861), .n5860(n5860), .n5859(n5859), .n5858(n5858), 
            .\REG.mem_55_15 (\REG.mem_55_15 ), .n5857(n5857), .\REG.mem_55_14 (\REG.mem_55_14 ), 
            .n5856(n5856), .n5855(n5855), .n5854(n5854), .\REG.mem_55_11 (\REG.mem_55_11 ), 
            .n5853(n5853), .\rd_sig_diff0_w[0] (rd_sig_diff0_w[0]), .n5852(n5852), 
            .n5851(n5851), .\REG.mem_55_8 (\REG.mem_55_8 ), .n5850(n5850), 
            .n5849(n5849), .\REG.mem_55_6 (\REG.mem_55_6 ), .n5848(n5848), 
            .\REG.mem_55_5 (\REG.mem_55_5 ), .n5847(n5847), .\REG.mem_55_4 (\REG.mem_55_4 ), 
            .n5846(n5846), .\REG.mem_55_3 (\REG.mem_55_3 ), .n5845(n5845), 
            .\REG.mem_55_2 (\REG.mem_55_2 ), .n5844(n5844), .\REG.mem_55_1 (\REG.mem_55_1 ), 
            .n5843(n5843), .\REG.mem_55_0 (\REG.mem_55_0 ), .n5842(n5842), 
            .n5841(n5841), .n5839(n5839), .n5838(n5838), .n5837(n5837), 
            .\REG.mem_16_15 (\REG.mem_16_15 ), .\REG.mem_18_15 (\REG.mem_18_15 ), 
            .\REG.mem_23_15 (\REG.mem_23_15 ), .n5836(n5836), .\REG.mem_25_4 (\REG.mem_25_4 ), 
            .\REG.mem_35_2 (\REG.mem_35_2 ), .\REG.mem_31_4 (\REG.mem_31_4 ), 
            .\REG.mem_38_2 (\REG.mem_38_2 ), .\REG.mem_39_2 (\REG.mem_39_2 ), 
            .\REG.mem_36_2 (\REG.mem_36_2 ), .\REG.mem_37_2 (\REG.mem_37_2 ), 
            .\REG.mem_10_15 (\REG.mem_10_15 ), .\REG.mem_11_15 (\REG.mem_11_15 ), 
            .\REG.mem_48_2 (\REG.mem_48_2 ), .\REG.mem_50_2 (\REG.mem_50_2 ), 
            .\REG.mem_8_4 (\REG.mem_8_4 ), .\REG.mem_9_4 (\REG.mem_9_4 ), 
            .\REG.mem_10_4 (\REG.mem_10_4 ), .\REG.mem_11_4 (\REG.mem_11_4 ), 
            .n5771(n5771), .\REG.mem_50_15 (\REG.mem_50_15 ), .n5770(n5770), 
            .\REG.mem_50_14 (\REG.mem_50_14 ), .n5769(n5769), .\REG.mem_50_13 (\REG.mem_50_13 ), 
            .n5768(n5768), .n5767(n5767), .\REG.mem_50_11 (\REG.mem_50_11 ), 
            .n5766(n5766), .n5765(n5765), .n5764(n5764), .\REG.mem_50_8 (\REG.mem_50_8 ), 
            .n5763(n5763), .n5762(n5762), .\REG.mem_50_6 (\REG.mem_50_6 ), 
            .n5761(n5761), .\REG.mem_50_5 (\REG.mem_50_5 ), .n5760(n5760), 
            .\REG.mem_50_4 (\REG.mem_50_4 ), .n5759(n5759), .n5758(n5758), 
            .n5757(n5757), .\REG.mem_14_4 (\REG.mem_14_4 ), .\REG.mem_15_4 (\REG.mem_15_4 ), 
            .n10873(n10873), .\REG.mem_12_4 (\REG.mem_12_4 ), .\REG.mem_13_4 (\REG.mem_13_4 ), 
            .n10582(n10582), .\fifo_data_out[14] (fifo_data_out[14]), .n10588(n10588), 
            .\fifo_data_out[15] (fifo_data_out[15]), .n5753(n5753), .\REG.mem_50_0 (\REG.mem_50_0 ), 
            .\REG.mem_3_14 (\REG.mem_3_14 ), .\REG.mem_6_14 (\REG.mem_6_14 ), 
            .\REG.mem_7_14 (\REG.mem_7_14 ), .\REG.mem_4_14 (\REG.mem_4_14 ), 
            .\REG.mem_5_14 (\REG.mem_5_14 ), .n5736(n5736), .\REG.mem_48_15 (\REG.mem_48_15 ), 
            .n5735(n5735), .\REG.mem_48_14 (\REG.mem_48_14 ), .n5734(n5734), 
            .\REG.mem_48_13 (\REG.mem_48_13 ), .n5733(n5733), .n5732(n5732), 
            .\REG.mem_48_11 (\REG.mem_48_11 ), .n5731(n5731), .n5730(n5730), 
            .n5729(n5729), .\REG.mem_48_8 (\REG.mem_48_8 ), .n5728(n5728), 
            .n5727(n5727), .\REG.mem_48_6 (\REG.mem_48_6 ), .n5726(n5726), 
            .\REG.mem_48_5 (\REG.mem_48_5 ), .n5725(n5725), .\REG.mem_48_4 (\REG.mem_48_4 ), 
            .n5724(n5724), .n10877(n10877), .\REG.mem_9_15 (\REG.mem_9_15 ), 
            .\REG.mem_8_15 (\REG.mem_8_15 ), .\REG.mem_31_7 (\REG.mem_31_7 ), 
            .n5723(n5723), .n5722(n5722), .n5721(n5721), .\REG.mem_48_0 (\REG.mem_48_0 ), 
            .n5720(n5720), .\REG.mem_47_15 (\REG.mem_47_15 ), .n5719(n5719), 
            .n5718(n5718), .\REG.mem_47_13 (\REG.mem_47_13 ), .n5717(n5717), 
            .\REG.mem_47_12 (\REG.mem_47_12 ), .n5716(n5716), .\REG.mem_47_11 (\REG.mem_47_11 ), 
            .n5715(n5715), .\REG.mem_47_10 (\REG.mem_47_10 ), .n5714(n5714), 
            .\REG.mem_47_9 (\REG.mem_47_9 ), .n5713(n5713), .n5712(n5712), 
            .\REG.mem_47_7 (\REG.mem_47_7 ), .n5711(n5711), .\REG.mem_47_6 (\REG.mem_47_6 ), 
            .n5710(n5710), .\REG.mem_47_5 (\REG.mem_47_5 ), .n5709(n5709), 
            .n5708(n5708), .n5707(n5707), .\REG.mem_47_2 (\REG.mem_47_2 ), 
            .n5706(n5706), .n5705(n5705), .\REG.mem_47_0 (\REG.mem_47_0 ), 
            .n5704(n5704), .\REG.mem_46_15 (\REG.mem_46_15 ), .n5703(n5703), 
            .\REG.mem_31_12 (\REG.mem_31_12 ), .n5702(n5702), .\REG.mem_46_13 (\REG.mem_46_13 ), 
            .n5701(n5701), .\REG.mem_46_12 (\REG.mem_46_12 ), .n5700(n5700), 
            .\REG.mem_46_11 (\REG.mem_46_11 ), .n5699(n5699), .\REG.mem_46_10 (\REG.mem_46_10 ), 
            .n5698(n5698), .\REG.mem_46_9 (\REG.mem_46_9 ), .n5697(n5697), 
            .n5696(n5696), .\REG.mem_46_7 (\REG.mem_46_7 ), .n5695(n5695), 
            .\REG.mem_46_6 (\REG.mem_46_6 ), .n5694(n5694), .\REG.mem_46_5 (\REG.mem_46_5 ), 
            .n5693(n5693), .n5692(n5692), .n5691(n5691), .\REG.mem_46_2 (\REG.mem_46_2 ), 
            .n5690(n5690), .n5689(n5689), .\REG.mem_46_0 (\REG.mem_46_0 ), 
            .n5688(n5688), .\REG.mem_45_15 (\REG.mem_45_15 ), .n5687(n5687), 
            .n5686(n5686), .\REG.mem_45_13 (\REG.mem_45_13 ), .n5685(n5685), 
            .\REG.mem_45_12 (\REG.mem_45_12 ), .n5684(n5684), .\REG.mem_45_11 (\REG.mem_45_11 ), 
            .n5683(n5683), .\REG.mem_45_10 (\REG.mem_45_10 ), .n5682(n5682), 
            .\REG.mem_45_9 (\REG.mem_45_9 ), .n5681(n5681), .n5680(n5680), 
            .\REG.mem_45_7 (\REG.mem_45_7 ), .n5679(n5679), .\REG.mem_45_6 (\REG.mem_45_6 ), 
            .n5678(n5678), .\REG.mem_45_5 (\REG.mem_45_5 ), .\REG.mem_38_6 (\REG.mem_38_6 ), 
            .\REG.mem_39_6 (\REG.mem_39_6 ), .\REG.mem_37_6 (\REG.mem_37_6 ), 
            .\REG.mem_36_6 (\REG.mem_36_6 ), .n5677(n5677), .\REG.mem_31_11 (\REG.mem_31_11 ), 
            .n5676(n5676), .\REG.mem_42_5 (\REG.mem_42_5 ), .\REG.mem_43_5 (\REG.mem_43_5 ), 
            .n5675(n5675), .\REG.mem_45_2 (\REG.mem_45_2 ), .n5674(n5674), 
            .n5673(n5673), .\REG.mem_45_0 (\REG.mem_45_0 ), .n5671(n5671), 
            .\REG.mem_44_15 (\REG.mem_44_15 ), .n5670(n5670), .n5669(n5669), 
            .\REG.mem_44_13 (\REG.mem_44_13 ), .n5668(n5668), .\REG.mem_44_12 (\REG.mem_44_12 ), 
            .n5666(n5666), .\REG.mem_44_11 (\REG.mem_44_11 ), .n5665(n5665), 
            .\REG.mem_44_10 (\REG.mem_44_10 ), .n5664(n5664), .\REG.mem_44_9 (\REG.mem_44_9 ), 
            .n5662(n5662), .n5661(n5661), .\REG.mem_44_7 (\REG.mem_44_7 ), 
            .n5660(n5660), .\REG.mem_44_6 (\REG.mem_44_6 ), .n5659(n5659), 
            .\REG.mem_44_5 (\REG.mem_44_5 ), .n5658(n5658), .n5657(n5657), 
            .n5656(n5656), .\REG.mem_44_2 (\REG.mem_44_2 ), .n5655(n5655), 
            .n5654(n5654), .\REG.mem_44_0 (\REG.mem_44_0 ), .n5653(n5653), 
            .\REG.mem_43_15 (\REG.mem_43_15 ), .n5652(n5652), .n5651(n5651), 
            .\REG.mem_43_13 (\REG.mem_43_13 ), .n5650(n5650), .\REG.mem_43_12 (\REG.mem_43_12 ), 
            .n5649(n5649), .\REG.mem_43_11 (\REG.mem_43_11 ), .n5648(n5648), 
            .\REG.mem_43_10 (\REG.mem_43_10 ), .n5647(n5647), .\REG.mem_43_9 (\REG.mem_43_9 ), 
            .n5646(n5646), .n5645(n5645), .\REG.mem_43_7 (\REG.mem_43_7 ), 
            .n5644(n5644), .\REG.mem_43_6 (\REG.mem_43_6 ), .\REG.mem_41_5 (\REG.mem_41_5 ), 
            .\REG.mem_40_5 (\REG.mem_40_5 ), .\REG.mem_23_1 (\REG.mem_23_1 ), 
            .\rd_addr_p1_w[0] (rd_addr_p1_w[0]), .\REG.mem_35_11 (\REG.mem_35_11 ), 
            .n5643(n5643), .n5642(n5642), .n5641(n5641), .n5640(n5640), 
            .\REG.mem_43_2 (\REG.mem_43_2 ), .n5639(n5639), .\REG.mem_43_1 (\REG.mem_43_1 ), 
            .n5638(n5638), .n5637(n5637), .\REG.mem_42_15 (\REG.mem_42_15 ), 
            .n5636(n5636), .n5635(n5635), .\REG.mem_42_13 (\REG.mem_42_13 ), 
            .n5634(n5634), .\REG.mem_42_12 (\REG.mem_42_12 ), .n5633(n5633), 
            .\REG.mem_42_11 (\REG.mem_42_11 ), .n5632(n5632), .\REG.mem_42_10 (\REG.mem_42_10 ), 
            .n5631(n5631), .\REG.mem_42_9 (\REG.mem_42_9 ), .n5630(n5630), 
            .n5629(n5629), .\REG.mem_42_7 (\REG.mem_42_7 ), .n4916(n4916), 
            .\REG.mem_31_6 (\REG.mem_31_6 ), .\REG.mem_23_2 (\REG.mem_23_2 ), 
            .\REG.mem_38_11 (\REG.mem_38_11 ), .\REG.mem_39_11 (\REG.mem_39_11 ), 
            .\REG.mem_37_11 (\REG.mem_37_11 ), .\REG.mem_36_11 (\REG.mem_36_11 ), 
            .n5628(n5628), .\REG.mem_42_6 (\REG.mem_42_6 ), .n5627(n5627), 
            .n5626(n5626), .n5625(n5625), .n5624(n5624), .\REG.mem_42_2 (\REG.mem_42_2 ), 
            .n5623(n5623), .\REG.mem_42_1 (\REG.mem_42_1 ), .n5622(n5622), 
            .n5621(n5621), .\REG.mem_41_15 (\REG.mem_41_15 ), .n5620(n5620), 
            .n5619(n5619), .\REG.mem_41_13 (\REG.mem_41_13 ), .n5618(n5618), 
            .\REG.mem_41_12 (\REG.mem_41_12 ), .n5617(n5617), .\REG.mem_41_11 (\REG.mem_41_11 ), 
            .n5616(n5616), .\REG.mem_41_10 (\REG.mem_41_10 ), .n5615(n5615), 
            .\REG.mem_41_9 (\REG.mem_41_9 ), .n5614(n5614), .n5613(n5613), 
            .\REG.mem_41_7 (\REG.mem_41_7 ), .\REG.mem_3_2 (\REG.mem_3_2 ), 
            .n5612(n5612), .\REG.mem_41_6 (\REG.mem_41_6 ), .n5611(n5611), 
            .n5610(n5610), .n5609(n5609), .n5608(n5608), .\REG.mem_41_2 (\REG.mem_41_2 ), 
            .n5607(n5607), .\REG.mem_41_1 (\REG.mem_41_1 ), .n5606(n5606), 
            .n5605(n5605), .\REG.mem_40_15 (\REG.mem_40_15 ), .n5604(n5604), 
            .n5603(n5603), .\REG.mem_40_13 (\REG.mem_40_13 ), .n5602(n5602), 
            .\REG.mem_40_12 (\REG.mem_40_12 ), .n5601(n5601), .\REG.mem_40_11 (\REG.mem_40_11 ), 
            .n5600(n5600), .\REG.mem_40_10 (\REG.mem_40_10 ), .n5599(n5599), 
            .\REG.mem_40_9 (\REG.mem_40_9 ), .n5598(n5598), .n5597(n5597), 
            .\REG.mem_40_7 (\REG.mem_40_7 ), .\REG.mem_25_9 (\REG.mem_25_9 ), 
            .n4904(n4904), .n4903(n4903), .n4901(n4901), .n4899(n4899), 
            .n5596(n5596), .\REG.mem_40_6 (\REG.mem_40_6 ), .n5595(n5595), 
            .n5594(n5594), .n5593(n5593), .n5592(n5592), .\REG.mem_40_2 (\REG.mem_40_2 ), 
            .n5591(n5591), .\REG.mem_40_1 (\REG.mem_40_1 ), .n5590(n5590), 
            .n5589(n5589), .n5588(n5588), .\REG.mem_39_14 (\REG.mem_39_14 ), 
            .n5587(n5587), .n5586(n5586), .\REG.mem_39_12 (\REG.mem_39_12 ), 
            .n5585(n5585), .n5584(n5584), .\REG.mem_39_10 (\REG.mem_39_10 ), 
            .n5583(n5583), .\REG.mem_39_9 (\REG.mem_39_9 ), .n5582(n5582), 
            .n5581(n5581), .n4898(n4898), .\REG.mem_14_1 (\REG.mem_14_1 ), 
            .\REG.mem_15_1 (\REG.mem_15_1 ), .DEBUG_5_c(DEBUG_5_c), .\REG.mem_13_1 (\REG.mem_13_1 ), 
            .\REG.mem_12_1 (\REG.mem_12_1 ), .\REG.mem_3_3 (\REG.mem_3_3 ), 
            .n5580(n5580), .n5579(n5579), .n5578(n5578), .\REG.mem_39_4 (\REG.mem_39_4 ), 
            .n5577(n5577), .n5576(n5576), .n5575(n5575), .\REG.mem_39_1 (\REG.mem_39_1 ), 
            .n5573(n5573), .n5572(n5572), .n5571(n5571), .\REG.mem_38_14 (\REG.mem_38_14 ), 
            .n5570(n5570), .n5569(n5569), .\REG.mem_38_12 (\REG.mem_38_12 ), 
            .n5568(n5568), .n5567(n5567), .\REG.mem_38_10 (\REG.mem_38_10 ), 
            .n5566(n5566), .\REG.mem_38_9 (\REG.mem_38_9 ), .n5565(n5565), 
            .n5564(n5564), .n5563(n5563), .n5562(n5562), .n5561(n5561), 
            .\REG.mem_38_4 (\REG.mem_38_4 ), .n5560(n5560), .n5559(n5559), 
            .n5558(n5558), .\REG.mem_38_1 (\REG.mem_38_1 ), .n5556(n5556), 
            .n5555(n5555), .n5554(n5554), .\REG.mem_37_14 (\REG.mem_37_14 ), 
            .n5553(n5553), .n5552(n5552), .\REG.mem_37_12 (\REG.mem_37_12 ), 
            .n5551(n5551), .n5550(n5550), .\REG.mem_37_10 (\REG.mem_37_10 ), 
            .n5549(n5549), .\REG.mem_37_9 (\REG.mem_37_9 ), .\REG.mem_25_13 (\REG.mem_25_13 ), 
            .\REG.out_raw[15] (\REG.out_raw [15]), .\REG.out_raw[14] (\REG.out_raw [14]), 
            .\REG.out_raw[13] (\REG.out_raw [13]), .\REG.out_raw[12] (\REG.out_raw [12]), 
            .\REG.out_raw[11] (\REG.out_raw [11]), .n5548(n5548), .n5547(n5547), 
            .n5546(n5546), .n5545(n5545), .n5544(n5544), .\REG.mem_37_4 (\REG.mem_37_4 ), 
            .n5543(n5543), .n5542(n5542), .n5541(n5541), .\REG.mem_37_1 (\REG.mem_37_1 ), 
            .n5540(n5540), .\REG.out_raw[10] (\REG.out_raw [10]), .\REG.out_raw[9] (\REG.out_raw [9]), 
            .\REG.out_raw[8] (\REG.out_raw [8]), .\REG.out_raw[7] (\REG.out_raw [7]), 
            .\REG.out_raw[6] (\REG.out_raw [6]), .\REG.out_raw[5] (\REG.out_raw [5]), 
            .\REG.out_raw[4] (\REG.out_raw [4]), .\REG.out_raw[3] (\REG.out_raw [3]), 
            .\REG.out_raw[2] (\REG.out_raw [2]), .\REG.out_raw[1] (\REG.out_raw [1]), 
            .n5526(n5526), .n5525(n5525), .\REG.mem_36_14 (\REG.mem_36_14 ), 
            .n5524(n5524), .n5523(n5523), .\REG.mem_36_12 (\REG.mem_36_12 ), 
            .n5522(n5522), .n5521(n5521), .\REG.mem_36_10 (\REG.mem_36_10 ), 
            .n5520(n5520), .\REG.mem_36_9 (\REG.mem_36_9 ), .n5519(n5519), 
            .n5518(n5518), .n5517(n5517), .n5516(n5516), .\rd_sig_diff0_w[2] (rd_sig_diff0_w[2]), 
            .n5515(n5515), .\REG.mem_36_4 (\REG.mem_36_4 ), .n5514(n5514), 
            .n5513(n5513), .n5512(n5512), .\REG.mem_36_1 (\REG.mem_36_1 ), 
            .n5511(n5511), .n5507(n5507), .n5506(n5506), .\REG.mem_35_14 (\REG.mem_35_14 ), 
            .n5505(n5505), .n5504(n5504), .\REG.mem_35_12 (\REG.mem_35_12 ), 
            .n5503(n5503), .n5502(n5502), .\REG.mem_35_10 (\REG.mem_35_10 ), 
            .n5501(n5501), .\REG.mem_35_9 (\REG.mem_35_9 ), .n5500(n5500), 
            .\rd_sig_diff0_w[1] (rd_sig_diff0_w[1]), .n5499(n5499), .\REG.mem_35_7 (\REG.mem_35_7 ), 
            .n5498(n5498), .\REG.mem_35_6 (\REG.mem_35_6 ), .n5497(n5497), 
            .\REG.mem_35_5 (\REG.mem_35_5 ), .n5496(n5496), .\REG.mem_35_4 (\REG.mem_35_4 ), 
            .n5495(n5495), .n5494(n5494), .n5493(n5493), .\REG.mem_35_1 (\REG.mem_35_1 ), 
            .n5492(n5492), .\REG.mem_6_3 (\REG.mem_6_3 ), .\REG.mem_7_3 (\REG.mem_7_3 ), 
            .\REG.mem_5_3 (\REG.mem_5_3 ), .\REG.mem_4_3 (\REG.mem_4_3 ), 
            .n5441(n5441), .n5440(n5440), .\REG.mem_31_14 (\REG.mem_31_14 ), 
            .n5439(n5439), .n5438(n5438), .n5437(n5437), .\REG.mem_25_1 (\REG.mem_25_1 ), 
            .n5436(n5436), .\REG.mem_31_10 (\REG.mem_31_10 ), .n58(n58), 
            .n5435(n5435), .\REG.mem_31_9 (\REG.mem_31_9 ), .n5434(n5434), 
            .\REG.mem_31_8 (\REG.mem_31_8 ), .n5433(n5433), .n5432(n5432), 
            .n5431(n5431), .n5430(n5430), .n5429(n5429), .n5428(n5428), 
            .n5427(n5427), .\REG.mem_31_1 (\REG.mem_31_1 ), .n5426(n5426), 
            .n26(n26), .DEBUG_1_c_c(DEBUG_1_c_c), .write_to_dc32_fifo_latched_N_425(write_to_dc32_fifo_latched_N_425), 
            .n5345(n5345), .n5344(n5344), .\REG.mem_25_14 (\REG.mem_25_14 ), 
            .n5343(n5343), .n5342(n5342), .n5341(n5341), .n5340(n5340), 
            .\REG.mem_25_10 (\REG.mem_25_10 ), .n5339(n5339), .n5338(n5338), 
            .\REG.mem_25_8 (\REG.mem_25_8 ), .n5337(n5337), .n5336(n5336), 
            .n5335(n5335), .n5334(n5334), .n5333(n5333), .\REG.mem_25_3 (\REG.mem_25_3 ), 
            .n5332(n5332), .n5331(n5331), .n5330(n5330), .\REG.mem_25_0 (\REG.mem_25_0 ), 
            .\REG.mem_14_15 (\REG.mem_14_15 ), .\REG.mem_15_15 (\REG.mem_15_15 ), 
            .\REG.mem_6_13 (\REG.mem_6_13 ), .\REG.mem_7_13 (\REG.mem_7_13 ), 
            .n5306(n5306), .n5305(n5305), .\REG.mem_23_14 (\REG.mem_23_14 ), 
            .n5304(n5304), .\REG.mem_23_13 (\REG.mem_23_13 ), .n5303(n5303), 
            .n5302(n5302), .n5301(n5301), .\REG.mem_23_10 (\REG.mem_23_10 ), 
            .n5300(n5300), .\REG.mem_23_9 (\REG.mem_23_9 ), .n5299(n5299), 
            .n5298(n5298), .\REG.mem_23_7 (\REG.mem_23_7 ), .n5297(n5297), 
            .\REG.mem_23_6 (\REG.mem_23_6 ), .n5296(n5296), .\REG.mem_23_5 (\REG.mem_23_5 ), 
            .n5295(n5295), .\REG.mem_23_4 (\REG.mem_23_4 ), .n5294(n5294), 
            .\REG.mem_23_3 (\REG.mem_23_3 ), .n5293(n5293), .n5292(n5292), 
            .n5290(n5290), .\REG.mem_23_0 (\REG.mem_23_0 ), .\rd_grey_sync_r[5] (rd_grey_sync_r[5]), 
            .\REG.mem_5_13 (\REG.mem_5_13 ), .\REG.mem_4_13 (\REG.mem_4_13 ), 
            .\rd_grey_sync_r[4] (rd_grey_sync_r[4]), .\rd_grey_sync_r[3] (rd_grey_sync_r[3]), 
            .\rd_grey_sync_r[2] (rd_grey_sync_r[2]), .\rd_grey_sync_r[1] (rd_grey_sync_r[1]), 
            .\REG.mem_13_15 (\REG.mem_13_15 ), .\REG.mem_12_15 (\REG.mem_12_15 ), 
            .n51(n51), .n19(n19), .\wr_addr_nxt_c[1] (wr_addr_nxt_c[1]), 
            .\REG.mem_10_0 (\REG.mem_10_0 ), .\REG.mem_11_0 (\REG.mem_11_0 ), 
            .\REG.mem_10_3 (\REG.mem_10_3 ), .\REG.mem_11_3 (\REG.mem_11_3 ), 
            .n5224(n5224), .n5223(n5223), .\REG.mem_18_14 (\REG.mem_18_14 ), 
            .n5222(n5222), .\REG.mem_18_13 (\REG.mem_18_13 ), .n5221(n5221), 
            .n5220(n5220), .\REG.mem_9_3 (\REG.mem_9_3 ), .\REG.mem_8_3 (\REG.mem_8_3 ), 
            .\REG.mem_9_0 (\REG.mem_9_0 ), .\REG.mem_8_0 (\REG.mem_8_0 ), 
            .\REG.mem_10_13 (\REG.mem_10_13 ), .\REG.mem_11_13 (\REG.mem_11_13 ), 
            .n52(n52), .\REG.mem_9_13 (\REG.mem_9_13 ), .\REG.mem_8_13 (\REG.mem_8_13 ), 
            .n20(n20), .n5219(n5219), .\REG.mem_18_10 (\REG.mem_18_10 ), 
            .n5218(n5218), .\REG.mem_18_9 (\REG.mem_18_9 ), .n5217(n5217), 
            .n5216(n5216), .n5215(n5215), .n5214(n5214), .\REG.mem_18_5 (\REG.mem_18_5 ), 
            .n5213(n5213), .\REG.mem_18_4 (\REG.mem_18_4 ), .n5212(n5212), 
            .\REG.mem_18_3 (\REG.mem_18_3 ), .n5211(n5211), .n5210(n5210), 
            .n5209(n5209), .\REG.mem_18_0 (\REG.mem_18_0 ), .\REG.mem_14_13 (\REG.mem_14_13 ), 
            .\REG.mem_15_13 (\REG.mem_15_13 ), .\REG.mem_13_13 (\REG.mem_13_13 ), 
            .\REG.mem_12_13 (\REG.mem_12_13 ), .\REG.mem_6_4 (\REG.mem_6_4 ), 
            .\REG.mem_7_4 (\REG.mem_7_4 ), .\REG.mem_5_4 (\REG.mem_5_4 ), 
            .\REG.mem_4_4 (\REG.mem_4_4 ), .get_next_word(get_next_word), 
            .n5188(n5188), .n5186(n5186), .\REG.mem_16_14 (\REG.mem_16_14 ), 
            .n5185(n5185), .\REG.mem_16_13 (\REG.mem_16_13 ), .\REG.mem_6_8 (\REG.mem_6_8 ), 
            .\REG.mem_7_8 (\REG.mem_7_8 ), .\REG.mem_3_6 (\REG.mem_3_6 ), 
            .n5184(n5184), .\REG.mem_5_8 (\REG.mem_5_8 ), .\REG.mem_4_8 (\REG.mem_4_8 ), 
            .\REG.mem_6_2 (\REG.mem_6_2 ), .\REG.mem_7_2 (\REG.mem_7_2 ), 
            .\REG.mem_5_2 (\REG.mem_5_2 ), .\REG.mem_4_2 (\REG.mem_4_2 ), 
            .rd_fifo_en_w(rd_fifo_en_w), .n5183(n5183), .n5182(n5182), 
            .\REG.mem_16_10 (\REG.mem_16_10 ), .n5181(n5181), .\REG.mem_16_9 (\REG.mem_16_9 ), 
            .n5180(n5180), .n5179(n5179), .n5178(n5178), .n5177(n5177), 
            .\REG.mem_16_5 (\REG.mem_16_5 ), .n5176(n5176), .\REG.mem_16_4 (\REG.mem_16_4 ), 
            .\REG.mem_3_12 (\REG.mem_3_12 ), .n5175(n5175), .\REG.mem_16_3 (\REG.mem_16_3 ), 
            .n5174(n5174), .n5173(n5173), .n5172(n5172), .\REG.mem_16_0 (\REG.mem_16_0 ), 
            .n5169(n5169), .n5168(n5168), .n5167(n5167), .n47(n47), 
            .n5166(n5166), .n15(n15_adj_60), .n5165(n5165), .n5164(n5164), 
            .\REG.mem_15_10 (\REG.mem_15_10 ), .n5163(n5163), .\REG.mem_15_9 (\REG.mem_15_9 ), 
            .n5162(n5162), .n5161(n5161), .n5160(n5160), .\REG.mem_15_6 (\REG.mem_15_6 ), 
            .n5159(n5159), .n5158(n5158), .n5157(n5157), .\REG.mem_15_3 (\REG.mem_15_3 ), 
            .n5156(n5156), .\REG.mem_15_2 (\REG.mem_15_2 ), .n5155(n5155), 
            .n5154(n5154), .\REG.mem_15_0 (\REG.mem_15_0 ), .n5153(n5153), 
            .n5152(n5152), .\REG.mem_6_6 (\REG.mem_6_6 ), .\REG.mem_7_6 (\REG.mem_7_6 ), 
            .n5151(n5151), .n5150(n5150), .n5149(n5149), .n5148(n5148), 
            .\REG.mem_14_10 (\REG.mem_14_10 ), .n5147(n5147), .\REG.mem_14_9 (\REG.mem_14_9 ), 
            .n5146(n5146), .n5145(n5145), .n5144(n5144), .\REG.mem_14_6 (\REG.mem_14_6 ), 
            .\REG.mem_4_6 (\REG.mem_4_6 ), .\REG.mem_5_6 (\REG.mem_5_6 ), 
            .n5143(n5143), .n5142(n5142), .n5141(n5141), .\REG.mem_14_3 (\REG.mem_14_3 ), 
            .n5140(n5140), .\REG.mem_14_2 (\REG.mem_14_2 ), .n5139(n5139), 
            .n5138(n5138), .\REG.mem_14_0 (\REG.mem_14_0 ), .n5137(n5137), 
            .n5136(n5136), .n5135(n5135), .n5134(n5134), .n5133(n5133), 
            .n5132(n5132), .\REG.mem_13_10 (\REG.mem_13_10 ), .\REG.mem_13_9 (\REG.mem_13_9 ), 
            .\REG.mem_12_9 (\REG.mem_12_9 ), .n5131(n5131), .n5130(n5130), 
            .n5129(n5129), .n5128(n5128), .\REG.mem_13_6 (\REG.mem_13_6 ), 
            .n5127(n5127), .n5126(n5126), .n5125(n5125), .\REG.mem_13_3 (\REG.mem_13_3 ), 
            .n5124(n5124), .\REG.mem_13_2 (\REG.mem_13_2 ), .n5123(n5123), 
            .\REG.mem_10_8 (\REG.mem_10_8 ), .\REG.mem_11_8 (\REG.mem_11_8 ), 
            .n5122(n5122), .\REG.mem_13_0 (\REG.mem_13_0 ), .n5121(n5121), 
            .n5120(n5120), .n5119(n5119), .n5118(n5118), .\REG.mem_3_9 (\REG.mem_3_9 ), 
            .\REG.mem_9_8 (\REG.mem_9_8 ), .\REG.mem_8_8 (\REG.mem_8_8 ), 
            .n5117(n5117), .\REG.mem_8_6 (\REG.mem_8_6 ), .\REG.mem_9_6 (\REG.mem_9_6 ), 
            .n5116(n5116), .\REG.mem_12_10 (\REG.mem_12_10 ), .\REG.mem_10_6 (\REG.mem_10_6 ), 
            .\REG.mem_11_6 (\REG.mem_11_6 ), .n53(n53), .n21(n21), .n5115(n5115), 
            .n5114(n5114), .n5113(n5113), .n5112(n5112), .\REG.mem_12_6 (\REG.mem_12_6 ), 
            .n50(n50), .n5111(n5111), .n18(n18), .\REG.mem_6_12 (\REG.mem_6_12 ), 
            .\REG.mem_7_12 (\REG.mem_7_12 ), .n5110(n5110), .n5109(n5109), 
            .\REG.mem_12_3 (\REG.mem_12_3 ), .n5108(n5108), .\REG.mem_12_2 (\REG.mem_12_2 ), 
            .\REG.mem_4_12 (\REG.mem_4_12 ), .\REG.mem_5_12 (\REG.mem_5_12 ), 
            .\REG.mem_10_2 (\REG.mem_10_2 ), .\REG.mem_11_2 (\REG.mem_11_2 ), 
            .n5107(n5107), .\REG.mem_9_2 (\REG.mem_9_2 ), .\REG.mem_8_2 (\REG.mem_8_2 ), 
            .n54(n54), .n22(n22), .n5106(n5106), .\REG.mem_12_0 (\REG.mem_12_0 ), 
            .\rd_addr_nxt_c_6__N_498[3] (rd_addr_nxt_c_6__N_498[3]), .n5105(n5105), 
            .n5104(n5104), .n5103(n5103), .n5102(n5102), .\REG.mem_11_12 (\REG.mem_11_12 ), 
            .n5101(n5101), .n5100(n5100), .\REG.mem_11_10 (\REG.mem_11_10 ), 
            .n5099(n5099), .n5098(n5098), .n5097(n5097), .n5096(n5096), 
            .n5095(n5095), .\REG.mem_11_5 (\REG.mem_11_5 ), .n5094(n5094), 
            .n5093(n5093), .n5092(n5092), .n5091(n5091), .\REG.mem_11_1 (\REG.mem_11_1 ), 
            .n5090(n5090), .n5089(n5089), .n5088(n5088), .\rd_addr_nxt_c_6__N_498[5] (rd_addr_nxt_c_6__N_498[5]), 
            .n5087(n5087), .n5086(n5086), .\REG.mem_10_12 (\REG.mem_10_12 ), 
            .n5085(n5085), .n5084(n5084), .\REG.mem_10_10 (\REG.mem_10_10 ), 
            .n5083(n5083), .n5082(n5082), .n5081(n5081), .n5080(n5080), 
            .n5079(n5079), .\REG.mem_10_5 (\REG.mem_10_5 ), .\REG.mem_10_1 (\REG.mem_10_1 ), 
            .\REG.mem_9_1 (\REG.mem_9_1 ), .\REG.mem_8_1 (\REG.mem_8_1 ), 
            .\rd_addr_nxt_c_6__N_498[2] (rd_addr_nxt_c_6__N_498[2]), .n56(n56), 
            .n24(n24_adj_61), .n5078(n5078), .n55(n55), .n23(n23), .n5077(n5077), 
            .n40(n40), .n8(n8_adj_59), .n5076(n5076), .n5075(n5075), 
            .n5074(n5074), .n5073(n5073), .n5072(n5072), .n5071(n5071), 
            .n5070(n5070), .\REG.mem_9_12 (\REG.mem_9_12 ), .n5069(n5069), 
            .n5068(n5068), .\REG.mem_9_10 (\REG.mem_9_10 ), .n5067(n5067), 
            .n5066(n5066), .n5065(n5065), .n57(n57), .n5064(n5064), 
            .n25(n25), .n5063(n5063), .\REG.mem_9_5 (\REG.mem_9_5 ), .n5062(n5062), 
            .n5061(n5061), .n5060(n5060), .n5059(n5059), .n5057(n5057), 
            .n5056(n5056), .n5055(n5055), .n5054(n5054), .n5053(n5053), 
            .\REG.mem_8_12 (\REG.mem_8_12 ), .n5052(n5052), .n5051(n5051), 
            .\REG.mem_8_10 (\REG.mem_8_10 ), .n5050(n5050), .n5049(n5049), 
            .n5048(n5048), .n5047(n5047), .n5046(n5046), .\REG.mem_8_5 (\REG.mem_8_5 ), 
            .n5045(n5045), .n5044(n5044), .n5043(n5043), .n5042(n5042), 
            .n5041(n5041), .n5040(n5040), .n5039(n5039), .n5038(n5038), 
            .n5037(n5037), .n5036(n5036), .n5035(n5035), .\REG.mem_7_10 (\REG.mem_7_10 ), 
            .n5034(n5034), .n5033(n5033), .n5032(n5032), .\REG.mem_7_7 (\REG.mem_7_7 ), 
            .n5031(n5031), .n5030(n5030), .\REG.mem_7_5 (\REG.mem_7_5 ), 
            .n5029(n5029), .n5028(n5028), .n5027(n5027), .n5026(n5026), 
            .n5025(n5025), .\REG.mem_7_0 (\REG.mem_7_0 ), .n5024(n5024), 
            .n5023(n5023), .n5022(n5022), .n5021(n5021), .n5020(n5020), 
            .n5019(n5019), .\REG.mem_6_10 (\REG.mem_6_10 ), .n5018(n5018), 
            .n5017(n5017), .n5016(n5016), .\REG.mem_6_7 (\REG.mem_6_7 ), 
            .n5015(n5015), .n5014(n5014), .\REG.mem_6_5 (\REG.mem_6_5 ), 
            .n5013(n5013), .n5012(n5012), .n5011(n5011), .n5010(n5010), 
            .n5009(n5009), .\REG.mem_6_0 (\REG.mem_6_0 ), .n5008(n5008), 
            .n5007(n5007), .n5006(n5006), .n5005(n5005), .n5004(n5004), 
            .n5003(n5003), .\REG.mem_5_10 (\REG.mem_5_10 ), .n5002(n5002), 
            .n5001(n5001), .n5000(n5000), .\REG.mem_5_7 (\REG.mem_5_7 ), 
            .n4999(n4999), .n4998(n4998), .\REG.mem_5_5 (\REG.mem_5_5 ), 
            .n4997(n4997), .n4996(n4996), .n4995(n4995), .n4994(n4994), 
            .n4993(n4993), .\REG.mem_5_0 (\REG.mem_5_0 ), .n4992(n4992), 
            .n4991(n4991), .n4990(n4990), .n4989(n4989), .n4988(n4988), 
            .n4987(n4987), .\REG.mem_4_10 (\REG.mem_4_10 ), .n4986(n4986), 
            .n4985(n4985), .n4984(n4984), .\REG.mem_4_7 (\REG.mem_4_7 ), 
            .n4983(n4983), .n4982(n4982), .\REG.mem_4_5 (\REG.mem_4_5 ), 
            .n4981(n4981), .n4980(n4980), .n4979(n4979), .n4978(n4978), 
            .n4977(n4977), .\REG.mem_4_0 (\REG.mem_4_0 ), .n4976(n4976), 
            .n4975(n4975), .n4974(n4974), .n4973(n4973), .n4972(n4972), 
            .n4971(n4971), .\REG.mem_3_10 (\REG.mem_3_10 ), .n4970(n4970), 
            .n4969(n4969), .\REG.mem_3_8 (\REG.mem_3_8 ), .FT_OE_N_420(FT_OE_N_420), 
            .n49(n49), .n17(n17), .n42(n42), .n10(n10), .n4968(n4968), 
            .\REG.mem_3_7 (\REG.mem_3_7 ), .n4967(n4967), .n4966(n4966), 
            .\REG.mem_3_5 (\REG.mem_3_5 ), .n4965(n4965), .n34(n34), .n4964(n4964), 
            .n4963(n4963), .n2(n2), .n4962(n4962), .n4961(n4961), .\REG.mem_3_0 (\REG.mem_3_0 ), 
            .n59(n59), .n27(n27), .n60(n60), .n28(n28), .n61(n61), 
            .n29(n29)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(547[21] 562[2])
    SB_LUT4 i3723_3_lut (.I0(\REG.mem_12_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n53), .I3(GND_net), .O(n5106));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3722_3_lut (.I0(\REG.mem_11_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n54), .I3(GND_net), .O(n5105));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(reset_all_w), .I3(GND_net), .O(empty_o_N_1149));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i3721_3_lut (.I0(\REG.mem_11_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n54), .I3(GND_net), .O(n5104));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3720_3_lut (.I0(\REG.mem_11_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n54), .I3(GND_net), .O(n5103));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3719_3_lut (.I0(\REG.mem_11_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n54), .I3(GND_net), .O(n5102));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3718_3_lut (.I0(\REG.mem_11_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n54), .I3(GND_net), .O(n5101));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3717_3_lut (.I0(\REG.mem_11_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n54), .I3(GND_net), .O(n5100));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3716_3_lut (.I0(\REG.mem_11_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n54), .I3(GND_net), .O(n5099));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3715_3_lut (.I0(\REG.mem_11_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n54), .I3(GND_net), .O(n5098));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3477_3_lut (.I0(tx_data_byte[1]), .I1(pc_data_rx[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4860));   // src/top.v(1074[8] 1141[4])
    defparam i3477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3714_3_lut (.I0(\REG.mem_11_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n54), .I3(GND_net), .O(n5097));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3713_3_lut (.I0(\REG.mem_11_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n54), .I3(GND_net), .O(n5096));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3712_3_lut (.I0(\REG.mem_11_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n54), .I3(GND_net), .O(n5095));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3711_3_lut (.I0(\REG.mem_11_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n54), .I3(GND_net), .O(n5094));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3710_3_lut (.I0(\REG.mem_11_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n54), .I3(GND_net), .O(n5093));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3709_3_lut (.I0(\REG.mem_11_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n54), .I3(GND_net), .O(n5092));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3709_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3708_3_lut (.I0(\REG.mem_11_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n54), .I3(GND_net), .O(n5091));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3707_3_lut (.I0(\REG.mem_11_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n54), .I3(GND_net), .O(n5090));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3706_3_lut (.I0(\REG.mem_10_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n55), .I3(GND_net), .O(n5089));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i949_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(n63), 
            .I3(state[2]), .O(n2034));   // src/timing_controller.v(51[11:16])
    defparam i949_4_lut_4_lut.LUT_INIT = 16'h0806;
    SB_LUT4 i3476_3_lut (.I0(tx_data_byte[2]), .I1(pc_data_rx[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4859));   // src/top.v(1074[8] 1141[4])
    defparam i3476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3472_3_lut (.I0(tx_data_byte[3]), .I1(pc_data_rx[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4855));   // src/top.v(1074[8] 1141[4])
    defparam i3472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3705_3_lut (.I0(\REG.mem_10_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n55), .I3(GND_net), .O(n5088));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3704_3_lut (.I0(\REG.mem_10_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n55), .I3(GND_net), .O(n5087));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3703_3_lut (.I0(\REG.mem_10_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n55), .I3(GND_net), .O(n5086));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3702_3_lut (.I0(\REG.mem_10_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n55), .I3(GND_net), .O(n5085));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3701_3_lut (.I0(\REG.mem_10_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n55), .I3(GND_net), .O(n5084));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3700_3_lut (.I0(\REG.mem_10_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n55), .I3(GND_net), .O(n5083));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3699_3_lut (.I0(\REG.mem_10_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n55), .I3(GND_net), .O(n5082));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3698_3_lut (.I0(\REG.mem_10_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n55), .I3(GND_net), .O(n5081));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3697_3_lut (.I0(\REG.mem_10_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n55), .I3(GND_net), .O(n5080));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3462_3_lut (.I0(tx_data_byte[4]), .I1(pc_data_rx[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4845));   // src/top.v(1074[8] 1141[4])
    defparam i3462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3696_3_lut (.I0(\REG.mem_10_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n55), .I3(GND_net), .O(n5079));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3695_3_lut (.I0(\REG.mem_10_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n55), .I3(GND_net), .O(n5078));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3694_3_lut (.I0(\REG.mem_10_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n55), .I3(GND_net), .O(n5077));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3693_3_lut (.I0(\REG.mem_10_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n55), .I3(GND_net), .O(n5076));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3692_3_lut (.I0(\REG.mem_10_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n55), .I3(GND_net), .O(n5075));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3455_3_lut (.I0(rx_shift_reg[5]), .I1(rx_shift_reg[4]), .I2(n4312), 
            .I3(GND_net), .O(n4838));   // src/spi.v(76[8] 221[4])
    defparam i3455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3691_3_lut (.I0(\REG.mem_10_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n55), .I3(GND_net), .O(n5074));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3690_3_lut (.I0(\REG.mem_9_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n56), .I3(GND_net), .O(n5073));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3689_3_lut (.I0(\REG.mem_9_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n56), .I3(GND_net), .O(n5072));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3688_3_lut (.I0(\REG.mem_9_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n56), .I3(GND_net), .O(n5071));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3687_3_lut (.I0(\REG.mem_9_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n56), .I3(GND_net), .O(n5070));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3686_3_lut (.I0(\REG.mem_9_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n56), .I3(GND_net), .O(n5069));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3453_3_lut (.I0(rx_shift_reg[6]), .I1(rx_shift_reg[5]), .I2(n4312), 
            .I3(GND_net), .O(n4836));   // src/spi.v(76[8] 221[4])
    defparam i3453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3685_3_lut (.I0(\REG.mem_9_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n56), .I3(GND_net), .O(n5068));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3684_3_lut (.I0(\REG.mem_9_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n56), .I3(GND_net), .O(n5067));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3683_3_lut (.I0(\REG.mem_9_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n56), .I3(GND_net), .O(n5066));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3682_3_lut (.I0(\REG.mem_9_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n56), .I3(GND_net), .O(n5065));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3681_3_lut (.I0(\REG.mem_9_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n56), .I3(GND_net), .O(n5064));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3680_3_lut (.I0(\REG.mem_9_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n56), .I3(GND_net), .O(n5063));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3679_3_lut (.I0(\REG.mem_9_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n56), .I3(GND_net), .O(n5062));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3678_3_lut (.I0(\REG.mem_9_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n56), .I3(GND_net), .O(n5061));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3677_3_lut (.I0(\REG.mem_9_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n56), .I3(GND_net), .O(n5060));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3676_3_lut (.I0(\REG.mem_9_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n56), .I3(GND_net), .O(n5059));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3674_3_lut (.I0(\REG.mem_9_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n56), .I3(GND_net), .O(n5057));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3673_3_lut (.I0(\REG.mem_8_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n57), .I3(GND_net), .O(n5056));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3672_3_lut (.I0(\REG.mem_8_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n57), .I3(GND_net), .O(n5055));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3671_3_lut (.I0(\REG.mem_8_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n57), .I3(GND_net), .O(n5054));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3670_3_lut (.I0(\REG.mem_8_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n57), .I3(GND_net), .O(n5053));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3669_3_lut (.I0(\REG.mem_8_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n57), .I3(GND_net), .O(n5052));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3668_3_lut (.I0(\REG.mem_8_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n57), .I3(GND_net), .O(n5051));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3667_3_lut (.I0(\REG.mem_8_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n57), .I3(GND_net), .O(n5050));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3666_3_lut (.I0(\REG.mem_8_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n57), .I3(GND_net), .O(n5049));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3665_3_lut (.I0(\REG.mem_8_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n57), .I3(GND_net), .O(n5048));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3664_3_lut (.I0(\REG.mem_8_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n57), .I3(GND_net), .O(n5047));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3663_3_lut (.I0(\REG.mem_8_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n57), .I3(GND_net), .O(n5046));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3662_3_lut (.I0(\REG.mem_8_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n57), .I3(GND_net), .O(n5045));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3661_3_lut (.I0(\REG.mem_8_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n57), .I3(GND_net), .O(n5044));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3660_3_lut (.I0(\REG.mem_8_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n57), .I3(GND_net), .O(n5043));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3659_3_lut (.I0(\REG.mem_8_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n57), .I3(GND_net), .O(n5042));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3658_3_lut (.I0(\REG.mem_8_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n57), .I3(GND_net), .O(n5041));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3657_3_lut (.I0(\REG.mem_7_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n58), .I3(GND_net), .O(n5040));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3656_3_lut (.I0(\REG.mem_7_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n58), .I3(GND_net), .O(n5039));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3655_3_lut (.I0(\REG.mem_7_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n58), .I3(GND_net), .O(n5038));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3654_3_lut (.I0(\REG.mem_7_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n58), .I3(GND_net), .O(n5037));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3653_3_lut (.I0(\REG.mem_7_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n58), .I3(GND_net), .O(n5036));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3652_3_lut (.I0(\REG.mem_7_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n58), .I3(GND_net), .O(n5035));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3651_3_lut (.I0(\REG.mem_7_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n58), .I3(GND_net), .O(n5034));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3650_3_lut (.I0(\REG.mem_7_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n58), .I3(GND_net), .O(n5033));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3649_3_lut (.I0(\REG.mem_7_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n58), .I3(GND_net), .O(n5032));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3648_3_lut (.I0(\REG.mem_7_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n58), .I3(GND_net), .O(n5031));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3647_3_lut (.I0(\REG.mem_7_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n58), .I3(GND_net), .O(n5030));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3646_3_lut (.I0(\REG.mem_7_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n58), .I3(GND_net), .O(n5029));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3645_3_lut (.I0(\REG.mem_7_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n58), .I3(GND_net), .O(n5028));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3644_3_lut (.I0(\REG.mem_7_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n58), .I3(GND_net), .O(n5027));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3643_3_lut (.I0(\REG.mem_7_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n58), .I3(GND_net), .O(n5026));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3642_3_lut (.I0(\REG.mem_7_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n58), .I3(GND_net), .O(n5025));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3641_3_lut (.I0(\REG.mem_6_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n59), .I3(GND_net), .O(n5024));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3554_2_lut_3_lut (.I0(fifo_data_out[2]), .I1(bluejay_data_out_31__N_736), 
            .I2(bluejay_data_out_31__N_737), .I3(GND_net), .O(n4937));   // src/bluejay_data.v(126[8] 148[4])
    defparam i3554_2_lut_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i3640_3_lut (.I0(\REG.mem_6_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n59), .I3(GND_net), .O(n5023));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3639_3_lut (.I0(\REG.mem_6_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n59), .I3(GND_net), .O(n5022));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3638_3_lut (.I0(\REG.mem_6_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n59), .I3(GND_net), .O(n5021));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3637_3_lut (.I0(\REG.mem_6_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n59), .I3(GND_net), .O(n5020));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3636_3_lut (.I0(\REG.mem_6_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n59), .I3(GND_net), .O(n5019));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3635_3_lut (.I0(\REG.mem_6_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n59), .I3(GND_net), .O(n5018));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3634_3_lut (.I0(\REG.mem_6_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n59), .I3(GND_net), .O(n5017));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3633_3_lut (.I0(\REG.mem_6_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n59), .I3(GND_net), .O(n5016));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3632_3_lut (.I0(\REG.mem_6_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n59), .I3(GND_net), .O(n5015));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3631_3_lut (.I0(\REG.mem_6_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n59), .I3(GND_net), .O(n5014));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3630_3_lut (.I0(\REG.mem_6_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n59), .I3(GND_net), .O(n5013));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3629_3_lut (.I0(\REG.mem_6_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n59), .I3(GND_net), .O(n5012));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3628_3_lut (.I0(\REG.mem_6_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n59), .I3(GND_net), .O(n5011));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3627_3_lut (.I0(\REG.mem_6_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n59), .I3(GND_net), .O(n5010));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3626_3_lut (.I0(\REG.mem_6_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n59), .I3(GND_net), .O(n5009));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3625_3_lut (.I0(\REG.mem_5_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n60), .I3(GND_net), .O(n5008));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3553_2_lut_3_lut (.I0(fifo_data_out[1]), .I1(bluejay_data_out_31__N_736), 
            .I2(bluejay_data_out_31__N_737), .I3(GND_net), .O(n4936));   // src/bluejay_data.v(126[8] 148[4])
    defparam i3553_2_lut_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i3624_3_lut (.I0(\REG.mem_5_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n60), .I3(GND_net), .O(n5007));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3623_3_lut (.I0(\REG.mem_5_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n60), .I3(GND_net), .O(n5006));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3622_3_lut (.I0(\REG.mem_5_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n60), .I3(GND_net), .O(n5005));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3621_3_lut (.I0(\REG.mem_5_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n60), .I3(GND_net), .O(n5004));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3620_3_lut (.I0(\REG.mem_5_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n60), .I3(GND_net), .O(n5003));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3620_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3619_3_lut (.I0(\REG.mem_5_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n60), .I3(GND_net), .O(n5002));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3618_3_lut (.I0(\REG.mem_5_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n60), .I3(GND_net), .O(n5001));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3617_3_lut (.I0(\REG.mem_5_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n60), .I3(GND_net), .O(n5000));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3616_3_lut (.I0(\REG.mem_5_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n60), .I3(GND_net), .O(n4999));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3615_3_lut (.I0(\REG.mem_5_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n60), .I3(GND_net), .O(n4998));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3614_3_lut (.I0(\REG.mem_5_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n60), .I3(GND_net), .O(n4997));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3613_3_lut (.I0(\REG.mem_5_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n60), .I3(GND_net), .O(n4996));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3612_3_lut (.I0(\REG.mem_5_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n60), .I3(GND_net), .O(n4995));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3611_3_lut (.I0(\REG.mem_5_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n60), .I3(GND_net), .O(n4994));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3610_3_lut (.I0(\REG.mem_5_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n60), .I3(GND_net), .O(n4993));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3609_3_lut (.I0(\REG.mem_4_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n61), .I3(GND_net), .O(n4992));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(reset_clk_counter[2]), .I1(reset_all_w_N_61), 
            .I2(reset_clk_counter[0]), .I3(reset_clk_counter[1]), .O(n10295));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'haaa6;
    SB_LUT4 i3608_3_lut (.I0(\REG.mem_4_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n61), .I3(GND_net), .O(n4991));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3608_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3607_3_lut (.I0(\REG.mem_4_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n61), .I3(GND_net), .O(n4990));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3606_3_lut (.I0(\REG.mem_4_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n61), .I3(GND_net), .O(n4989));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3605_3_lut (.I0(\REG.mem_4_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n61), .I3(GND_net), .O(n4988));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3604_3_lut (.I0(\REG.mem_4_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n61), .I3(GND_net), .O(n4987));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3603_3_lut (.I0(\REG.mem_4_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n61), .I3(GND_net), .O(n4986));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3602_3_lut (.I0(\REG.mem_4_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n61), .I3(GND_net), .O(n4985));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3601_3_lut (.I0(\REG.mem_4_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n61), .I3(GND_net), .O(n4984));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3600_3_lut (.I0(\REG.mem_4_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n61), .I3(GND_net), .O(n4983));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3599_3_lut (.I0(\REG.mem_4_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n61), .I3(GND_net), .O(n4982));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3598_3_lut (.I0(\REG.mem_4_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n61), .I3(GND_net), .O(n4981));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3597_3_lut (.I0(\REG.mem_4_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n61), .I3(GND_net), .O(n4980));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3596_3_lut (.I0(\REG.mem_4_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n61), .I3(GND_net), .O(n4979));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3595_3_lut (.I0(\REG.mem_4_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n61), .I3(GND_net), .O(n4978));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3594_3_lut (.I0(\REG.mem_4_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n61), .I3(GND_net), .O(n4977));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3593_3_lut (.I0(\REG.mem_3_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n62), .I3(GND_net), .O(n4976));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3592_3_lut (.I0(\REG.mem_3_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n62), .I3(GND_net), .O(n4975));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3591_3_lut (.I0(\REG.mem_3_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n62), .I3(GND_net), .O(n4974));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3590_3_lut (.I0(\REG.mem_3_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n62), .I3(GND_net), .O(n4973));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3589_3_lut (.I0(\REG.mem_3_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n62), .I3(GND_net), .O(n4972));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3588_3_lut (.I0(\REG.mem_3_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n62), .I3(GND_net), .O(n4971));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3587_3_lut (.I0(\REG.mem_3_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n62), .I3(GND_net), .O(n4970));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3586_3_lut (.I0(\REG.mem_3_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n62), .I3(GND_net), .O(n4969));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8368_2_lut_3_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(reset_clk_counter[1]), .I3(GND_net), .O(n10064));   // src/top.v(259[27:51])
    defparam i8368_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i4729_2_lut_3_lut (.I0(fifo_data_out[0]), .I1(bluejay_data_out_31__N_736), 
            .I2(bluejay_data_out_31__N_737), .I3(GND_net), .O(n6112));   // src/bluejay_data.v(126[8] 148[4])
    defparam i4729_2_lut_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_2_lut_3_lut_adj_90 (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(reset_clk_counter[1]), .I3(GND_net), .O(n10291));   // src/top.v(259[27:51])
    defparam i1_2_lut_3_lut_adj_90.LUT_INIT = 16'hd2d2;
    SB_LUT4 i1_4_lut_4_lut (.I0(is_tx_fifo_full_flag), .I1(n10917), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4723_3_lut_4_lut (.I0(r_SM_Main_2__N_844[0]), .I1(fifo_read_cmd), 
            .I2(is_fifo_empty_flag), .I3(tx_uart_active_flag), .O(n6106));   // src/top.v(910[8] 928[4])
    defparam i4723_3_lut_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_95[1]), .I1(r_SM_Main_2__N_841[1]), 
            .I2(r_SM_Main_adj_95[0]), .I3(r_SM_Main_adj_95[2]), .O(n13865));   // src/uart_tx.v(38[10] 141[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i3533_2_lut_3_lut (.I0(reset_per_frame), .I1(DEBUG_3_c), .I2(get_next_word), 
            .I3(GND_net), .O(n4916));   // src/fifo_dc_32_lut_gen.v(751[29] 761[32])
    defparam i3533_2_lut_3_lut.LUT_INIT = 16'h1010;
    clock clock_inst (.GND_net(GND_net), .VCC_net(VCC_net), .ICE_SYSCLK_c(ICE_SYSCLK_c), 
          .pll_clk_unbuf(pll_clk_unbuf)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(222[7] 228[3])
    SB_LUT4 i1_2_lut_4_lut_adj_91 (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(wr_addr_r_adj_118[0]), .I3(rd_addr_r_adj_121[0]), .O(n4_adj_58));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_2_lut_4_lut_adj_91.LUT_INIT = 16'h0220;
    SB_LUT4 i3451_3_lut (.I0(rx_shift_reg[7]), .I1(rx_shift_reg[6]), .I2(n4312), 
            .I3(GND_net), .O(n4834));   // src/spi.v(76[8] 221[4])
    defparam i3451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10380_4_lut (.I0(tx_data_byte[0]), .I1(tx_data_byte[1]), .I2(tx_data_byte[6]), 
            .I3(n10983), .O(multi_byte_spi_trans_flag_r_N_72));   // src/top.v(1123[10:31])
    defparam i10380_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i9145_4_lut (.I0(tx_data_byte[3]), .I1(tx_data_byte[2]), .I2(tx_data_byte[4]), 
            .I3(n10913), .O(n10983));
    defparam i9145_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i9076_2_lut (.I0(tx_data_byte[5]), .I1(tx_data_byte[7]), .I2(GND_net), 
            .I3(GND_net), .O(n10913));
    defparam i9076_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3585_3_lut (.I0(\REG.mem_3_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n62), .I3(GND_net), .O(n4968));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3584_3_lut (.I0(\REG.mem_3_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n62), .I3(GND_net), .O(n4967));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3584_3_lut.LUT_INIT = 16'hcaca;
    \uart_rx(CLKS_PER_BIT=20)  pc_rx (.r_SM_Main({r_SM_Main}), .SLM_CLK_c(SLM_CLK_c), 
            .r_Rx_Data(r_Rx_Data), .GND_net(GND_net), .n4(n4), .n4_adj_1(n4_adj_78), 
            .n6105(n6105), .pc_data_rx({pc_data_rx}), .n10406(n10406), 
            .VCC_net(VCC_net), .debug_led3(debug_led3), .n7473(n7473), 
            .n6082(n6082), .n6081(n6081), .n6079(n6079), .n6078(n6078), 
            .n6077(n6077), .n6075(n6075), .n6074(n6074), .\r_SM_Main_2__N_765[2] (r_SM_Main_2__N_765[2]), 
            .n4_adj_2(n4_adj_77), .n10345(n10345), .UART_RX_c(UART_RX_c), 
            .n4248(n4248), .n4253(n4253)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(699[42] 704[3])
    SB_LUT4 i3583_3_lut (.I0(\REG.mem_3_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n62), .I3(GND_net), .O(n4966));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3582_3_lut (.I0(\REG.mem_3_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n62), .I3(GND_net), .O(n4965));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3581_3_lut (.I0(\REG.mem_3_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n62), .I3(GND_net), .O(n4964));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3441_3_lut (.I0(tx_data_byte[0]), .I1(pc_data_rx[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4824));   // src/top.v(1074[8] 1141[4])
    defparam i3441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3580_3_lut (.I0(\REG.mem_3_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n62), .I3(GND_net), .O(n4963));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3580_3_lut.LUT_INIT = 16'hcaca;
    FIFO_Quad_Word tx_fifo (.rd_fifo_en_w(rd_fifo_en_w_adj_56), .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r [7]), 
            .SLM_CLK_c(SLM_CLK_c), .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r [6]), 
            .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r [5]), .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r [0]), 
            .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r [4]), .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r [3]), 
            .rd_addr_r({rd_addr_r_adj_121}), .reset_all_w(reset_all_w), 
            .n8(n8), .wr_addr_r({wr_addr_r_adj_118}), .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r [2]), 
            .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r [1]), .GND_net(GND_net), 
            .\rd_addr_p1_w[2] (rd_addr_p1_w_adj_123[2]), .n14025(n14025), 
            .n6127(n6127), .VCC_net(VCC_net), .\fifo_temp_output[1] (fifo_temp_output[1]), 
            .n10430(n10430), .is_tx_fifo_full_flag(is_tx_fifo_full_flag), 
            .n6088(n6088), .\fifo_temp_output[0] (fifo_temp_output[0]), 
            .\wr_addr_p1_w[2] (wr_addr_p1_w_adj_120[2]), .n1(n1), .n10226(n10226), 
            .n5989(n5989), .n5311(n5311), .\fifo_temp_output[4] (fifo_temp_output[4]), 
            .n5314(n5314), .\fifo_temp_output[5] (fifo_temp_output[5]), 
            .rx_buf_byte({rx_buf_byte}), .n5868(n5868), .n4882(n4882), 
            .\fifo_temp_output[2] (fifo_temp_output[2]), .n4887(n4887), 
            .\fifo_temp_output[3] (fifo_temp_output[3]), .n5536(n5536), 
            .\fifo_temp_output[6] (fifo_temp_output[6]), .n5539(n5539), 
            .\fifo_temp_output[7] (fifo_temp_output[7]), .n10786(n10786), 
            .is_fifo_empty_flag(is_fifo_empty_flag), .n4919(n4919), .n4922(n4922), 
            .fifo_write_cmd(fifo_write_cmd), .wr_fifo_en_w(wr_fifo_en_w), 
            .n4878(n4878), .rd_fifo_en_prev_r(rd_fifo_en_prev_r), .fifo_read_cmd(fifo_read_cmd)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(933[16] 949[2])
    SB_LUT4 i3579_3_lut (.I0(\REG.mem_3_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n62), .I3(GND_net), .O(n4962));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3579_3_lut.LUT_INIT = 16'hcaca;
    spi spi0 (.\tx_data_byte[3] (tx_data_byte[3]), .n2086(n2086), .GND_net(GND_net), 
        .\tx_data_byte[4] (tx_data_byte[4]), .SEN_c_1(SEN_c_1), .SLM_CLK_c(SLM_CLK_c), 
        .\tx_data_byte[5] (tx_data_byte[5]), .SOUT_c(SOUT_c), .n4312(n4312), 
        .\rx_shift_reg[0] (rx_shift_reg[0]), .\tx_data_byte[6] (tx_data_byte[6]), 
        .n4319(n4319), .SDAT_c_15(SDAT_c_15), .\tx_data_byte[7] (tx_data_byte[7]), 
        .tx_addr_byte({tx_addr_byte}), .VCC_net(VCC_net), .n10428(n10428), 
        .\tx_shift_reg[0] (tx_shift_reg[0]), .n6060(n6060), .rx_buf_byte({rx_buf_byte}), 
        .n6059(n6059), .n6058(n6058), .n6057(n6057), .n6056(n6056), 
        .n6055(n6055), .n6054(n6054), .spi_rx_byte_ready(spi_rx_byte_ready), 
        .SCK_c_0(SCK_c_0), .spi_start_transfer_r(spi_start_transfer_r), 
        .n4897(n4897), .n4888(n4888), .\rx_shift_reg[1] (rx_shift_reg[1]), 
        .n4883(n4883), .\rx_shift_reg[2] (rx_shift_reg[2]), .n4877(n4877), 
        .\rx_shift_reg[3] (rx_shift_reg[3]), .n4869(n4869), .\rx_shift_reg[4] (rx_shift_reg[4]), 
        .n4838(n4838), .\rx_shift_reg[5] (rx_shift_reg[5]), .multi_byte_spi_trans_flag_r(multi_byte_spi_trans_flag_r), 
        .n4836(n4836), .\rx_shift_reg[6] (rx_shift_reg[6]), .n4834(n4834), 
        .\rx_shift_reg[7] (rx_shift_reg[7]), .\tx_data_byte[2] (tx_data_byte[2]), 
        .\tx_data_byte[1] (tx_data_byte[1]), .n3495(n3495)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(833[5] 857[2])
    SB_LUT4 i3578_3_lut (.I0(\REG.mem_3_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n62), .I3(GND_net), .O(n4961));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3578_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3518_2_lut_4_lut (.I0(reset_per_frame), .I1(rd_addr_r[0]), 
            .I2(rd_addr_p1_w[0]), .I3(rd_fifo_en_w), .O(n4901));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i3518_2_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i3536_4_lut_4_lut (.I0(reset_all_w), .I1(rd_addr_r_adj_121[1]), 
            .I2(rd_addr_r_adj_121[0]), .I3(rd_fifo_en_w_adj_56), .O(n4919));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i3536_4_lut_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i4153_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[6]), 
            .I2(\mem_LUT.data_raw_r [6]), .I3(n4459), .O(n5536));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4153_4_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4156_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[7]), 
            .I2(\mem_LUT.data_raw_r [7]), .I3(n4459), .O(n5539));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4156_4_lut_4_lut.LUT_INIT = 16'h5044;
    \uart_tx(CLKS_PER_BIT=20)  pc_tx (.UART_TX_c(UART_TX_c), .SLM_CLK_c(SLM_CLK_c), 
            .r_SM_Main({r_SM_Main_adj_95}), .GND_net(GND_net), .\r_SM_Main_2__N_841[1] (r_SM_Main_2__N_841[1]), 
            .\r_SM_Main_2__N_844[0] (r_SM_Main_2__N_844[0]), .n3794(n3794), 
            .VCC_net(VCC_net), .n13865(n13865), .n10805(n10805), .n4890(n4890), 
            .r_Tx_Data({r_Tx_Data}), .n4889(n4889), .tx_uart_active_flag(tx_uart_active_flag), 
            .n5192(n5192), .n5191(n5191), .n5190(n5190), .n5189(n5189), 
            .n5187(n5187), .n5171(n5171), .n5170(n5170)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(768[42] 777[3])
    usb3_if usb3_if_inst (.reset_per_frame(reset_per_frame), .reset_per_frame_latched(reset_per_frame_latched), 
            .SLM_CLK_c(SLM_CLK_c), .DEBUG_3_c(DEBUG_3_c), .DEBUG_2_c(DEBUG_2_c), 
            .FIFO_CLK_c(FIFO_CLK_c), .\dc32_fifo_data_in[0] (dc32_fifo_data_in[0]), 
            .DEBUG_5_c(DEBUG_5_c), .buffer_switch_done(buffer_switch_done), 
            .buffer_switch_done_latched(buffer_switch_done_latched), .VCC_net(VCC_net), 
            .FT_OE_c(FT_OE_c), .n571(n571), .GND_net(GND_net), .n575(n575), 
            .write_to_dc32_fifo_latched_N_425(write_to_dc32_fifo_latched_N_425), 
            .n2352(n2352), .n4911(n4911), .n4910(n4910), .n4907(n4907), 
            .FIFO_D15_c_15(FIFO_D15_c_15), .FIFO_D14_c_14(FIFO_D14_c_14), 
            .FIFO_D13_c_13(FIFO_D13_c_13), .FIFO_D12_c_12(FIFO_D12_c_12), 
            .FIFO_D11_c_11(FIFO_D11_c_11), .FIFO_D10_c_10(FIFO_D10_c_10), 
            .FIFO_D9_c_9(FIFO_D9_c_9), .FIFO_D8_c_8(FIFO_D8_c_8), .FIFO_D7_c_7(FIFO_D7_c_7), 
            .FIFO_D6_c_6(FIFO_D6_c_6), .FIFO_D5_c_5(FIFO_D5_c_5), .FIFO_D4_c_4(FIFO_D4_c_4), 
            .FIFO_D3_c_3(FIFO_D3_c_3), .FIFO_D2_c_2(FIFO_D2_c_2), .FIFO_D1_c_1(FIFO_D1_c_1), 
            .dc32_fifo_almost_full(dc32_fifo_almost_full), .\dc32_fifo_data_in[15] (dc32_fifo_data_in[15]), 
            .\dc32_fifo_data_in[14] (dc32_fifo_data_in[14]), .\dc32_fifo_data_in[13] (dc32_fifo_data_in[13]), 
            .\dc32_fifo_data_in[12] (dc32_fifo_data_in[12]), .\dc32_fifo_data_in[11] (dc32_fifo_data_in[11]), 
            .\dc32_fifo_data_in[10] (dc32_fifo_data_in[10]), .\dc32_fifo_data_in[9] (dc32_fifo_data_in[9]), 
            .\dc32_fifo_data_in[8] (dc32_fifo_data_in[8]), .\dc32_fifo_data_in[7] (dc32_fifo_data_in[7]), 
            .\dc32_fifo_data_in[6] (dc32_fifo_data_in[6]), .\dc32_fifo_data_in[5] (dc32_fifo_data_in[5]), 
            .\dc32_fifo_data_in[4] (dc32_fifo_data_in[4]), .\dc32_fifo_data_in[3] (dc32_fifo_data_in[3]), 
            .\dc32_fifo_data_in[2] (dc32_fifo_data_in[2]), .\dc32_fifo_data_in[1] (dc32_fifo_data_in[1]), 
            .DEBUG_1_c_c(DEBUG_1_c_c), .FT_OE_N_420(FT_OE_N_420)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(513[9] 530[3])
    
endmodule
//
// Verilog Description of module timing_controller
//

module timing_controller (state, SLM_CLK_c, n1879, GND_net, n10514, 
            VCC_net, n10808, reset_per_frame, n1774, n7386, INVERT_c_3, 
            buffer_switch_done, n4245, n7568, n7590, n4192, n63, 
            n10831, UPDATE_c_2) /* synthesis syn_module_defined=1 */ ;
    output [3:0]state;
    input SLM_CLK_c;
    input n1879;
    input GND_net;
    input n10514;
    input VCC_net;
    input n10808;
    output reset_per_frame;
    input n1774;
    input n7386;
    output INVERT_c_3;
    output buffer_switch_done;
    output n4245;
    output n7568;
    input n7590;
    output n4192;
    output n63;
    output n10831;
    output UPDATE_c_2;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n13875;
    wire [3:0]state_3__N_80;
    
    wire n10833, n10814, n1951;
    wire [31:0]n1880;
    wire [31:0]n1952;
    wire [31:0]n506;
    
    wire n4491;
    wire [31:0]state_timeout_counter;   // src/timing_controller.v(52[12:33])
    
    wire n4809, n12053, n12051, n10121, n10122, n10105, n10106, 
        n12050, n10104, n12043, n10120, n10103, n12044, n10119, 
        n10102, n10118, n12036, n10117, n10132, n10131, n12045, 
        n10116, n12046, n10115, n10130, n10114, n12047, n10113, 
        n10129, n10128, n10127, n10112, n12048, n10111, n10126, 
        n12049, n10110, n10109, n12039, n10125, n12040, n10124, 
        n12041, n10123, n10108;
    wire [3:0]n968;
    
    wire n10107, n4806, n12054, n10823, n12042, n12106, n2033, 
        n4496, n10837, n38, n52, n56, n54, n55, n53, n50, 
        n58, n62, n49, n7570, n7, n12202, n5;
    
    SB_LUT4 i3_4_lut (.I0(state[3]), .I1(state[0]), .I2(state[1]), .I3(state[2]), 
            .O(n13875));
    defparam i3_4_lut.LUT_INIT = 16'h0400;
    SB_DFFE state_i0 (.Q(state[0]), .C(SLM_CLK_c), .E(n10833), .D(state_3__N_80[0]));   // src/timing_controller.v(56[8] 132[4])
    SB_LUT4 mux_898_i25_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[24]), .O(n1952[24]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i25_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i24_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[23]), .O(n1952[23]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i24_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i23_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[22]), .O(n1952[22]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i23_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i21_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[20]), .O(n1952[20]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i21_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i20_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[19]), .O(n1952[19]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i20_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i19_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[18]), .O(n1952[18]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i19_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i16_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[15]), .O(n1952[15]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i16_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i15_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[14]), .O(n1952[14]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i15_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i13_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[12]), .O(n1952[12]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i13_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i10_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[9]), .O(n1952[9]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i10_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i11_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[10]), .O(n1952[10]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i11_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i4_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[3]), .O(n1952[3]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i4_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_DFFESR state_timeout_counter_i0_i31 (.Q(state_timeout_counter[31]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[31]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i30 (.Q(state_timeout_counter[30]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[30]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_LUT4 mux_890_i2_3_lut (.I0(n12053), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[1]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i2_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i3_3_lut (.I0(n12051), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[2]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFE state_i3 (.Q(state[3]), .C(SLM_CLK_c), .E(VCC_net), .D(n10514));   // src/timing_controller.v(56[8] 132[4])
    SB_DFF invert_55_i0 (.Q(reset_per_frame), .C(SLM_CLK_c), .D(n10808));   // src/timing_controller.v(62[5] 131[12])
    SB_DFFESR state_timeout_counter_i0_i29 (.Q(state_timeout_counter[29]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[29]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i28 (.Q(state_timeout_counter[28]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[28]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i27 (.Q(state_timeout_counter[27]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[27]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i26 (.Q(state_timeout_counter[26]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[26]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i25 (.Q(state_timeout_counter[25]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[25]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i21 (.Q(state_timeout_counter[21]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[21]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i17 (.Q(state_timeout_counter[17]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[17]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i16 (.Q(state_timeout_counter[16]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[16]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i13 (.Q(state_timeout_counter[13]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[13]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i11 (.Q(state_timeout_counter[11]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[11]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_CARRY sub_31_add_2_22 (.CI(n10121), .I0(state_timeout_counter[20]), 
            .I1(VCC_net), .CO(n10122));
    SB_CARRY sub_31_add_2_6 (.CI(n10105), .I0(state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n10106));
    SB_LUT4 sub_31_add_2_5_lut (.I0(n1774), .I1(state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n10104), .O(n12050)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_21_lut (.I0(n1774), .I1(state_timeout_counter[19]), 
            .I2(VCC_net), .I3(n10120), .O(n12043)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_21 (.CI(n10120), .I0(state_timeout_counter[19]), 
            .I1(VCC_net), .CO(n10121));
    SB_CARRY sub_31_add_2_5 (.CI(n10104), .I0(state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n10105));
    SB_LUT4 sub_31_add_2_4_lut (.I0(n7386), .I1(state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n10103), .O(n12051)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_31_add_2_20_lut (.I0(n1774), .I1(state_timeout_counter[18]), 
            .I2(VCC_net), .I3(n10119), .O(n12044)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_20 (.CI(n10119), .I0(state_timeout_counter[18]), 
            .I1(VCC_net), .CO(n10120));
    SB_CARRY sub_31_add_2_4 (.CI(n10103), .I0(state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n10104));
    SB_LUT4 sub_31_add_2_3_lut (.I0(n1774), .I1(state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n10102), .O(n12053)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_19_lut (.I0(GND_net), .I1(state_timeout_counter[17]), 
            .I2(VCC_net), .I3(n10118), .O(n506[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_19 (.CI(n10118), .I0(state_timeout_counter[17]), 
            .I1(VCC_net), .CO(n10119));
    SB_CARRY sub_31_add_2_3 (.CI(n10102), .I0(state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n10103));
    SB_LUT4 sub_31_add_2_2_lut (.I0(n7386), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n12036)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_31_add_2_18_lut (.I0(GND_net), .I1(state_timeout_counter[16]), 
            .I2(VCC_net), .I3(n10117), .O(n506[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_33_lut (.I0(GND_net), .I1(state_timeout_counter[31]), 
            .I2(VCC_net), .I3(n10132), .O(n506[31])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_32_lut (.I0(GND_net), .I1(state_timeout_counter[30]), 
            .I2(VCC_net), .I3(n10131), .O(n506[30])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_18 (.CI(n10117), .I0(state_timeout_counter[16]), 
            .I1(VCC_net), .CO(n10118));
    SB_CARRY sub_31_add_2_2 (.CI(VCC_net), .I0(state_timeout_counter[0]), 
            .I1(GND_net), .CO(n10102));
    SB_LUT4 sub_31_add_2_17_lut (.I0(n1774), .I1(state_timeout_counter[15]), 
            .I2(VCC_net), .I3(n10116), .O(n12045)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_32 (.CI(n10131), .I0(state_timeout_counter[30]), 
            .I1(VCC_net), .CO(n10132));
    SB_CARRY sub_31_add_2_17 (.CI(n10116), .I0(state_timeout_counter[15]), 
            .I1(VCC_net), .CO(n10117));
    SB_LUT4 sub_31_add_2_16_lut (.I0(n1774), .I1(state_timeout_counter[14]), 
            .I2(VCC_net), .I3(n10115), .O(n12046)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_31_lut (.I0(GND_net), .I1(state_timeout_counter[29]), 
            .I2(VCC_net), .I3(n10130), .O(n506[29])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_16 (.CI(n10115), .I0(state_timeout_counter[14]), 
            .I1(VCC_net), .CO(n10116));
    SB_LUT4 sub_31_add_2_15_lut (.I0(GND_net), .I1(state_timeout_counter[13]), 
            .I2(VCC_net), .I3(n10114), .O(n506[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_31 (.CI(n10130), .I0(state_timeout_counter[29]), 
            .I1(VCC_net), .CO(n10131));
    SB_CARRY sub_31_add_2_15 (.CI(n10114), .I0(state_timeout_counter[13]), 
            .I1(VCC_net), .CO(n10115));
    SB_LUT4 sub_31_add_2_14_lut (.I0(n1774), .I1(state_timeout_counter[12]), 
            .I2(VCC_net), .I3(n10113), .O(n12047)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_30_lut (.I0(GND_net), .I1(state_timeout_counter[28]), 
            .I2(VCC_net), .I3(n10129), .O(n506[28])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_30 (.CI(n10129), .I0(state_timeout_counter[28]), 
            .I1(VCC_net), .CO(n10130));
    SB_LUT4 sub_31_add_2_29_lut (.I0(GND_net), .I1(state_timeout_counter[27]), 
            .I2(VCC_net), .I3(n10128), .O(n506[27])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_29 (.CI(n10128), .I0(state_timeout_counter[27]), 
            .I1(VCC_net), .CO(n10129));
    SB_LUT4 sub_31_add_2_28_lut (.I0(GND_net), .I1(state_timeout_counter[26]), 
            .I2(VCC_net), .I3(n10127), .O(n506[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_14 (.CI(n10113), .I0(state_timeout_counter[12]), 
            .I1(VCC_net), .CO(n10114));
    SB_LUT4 sub_31_add_2_13_lut (.I0(GND_net), .I1(state_timeout_counter[11]), 
            .I2(VCC_net), .I3(n10112), .O(n506[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_28 (.CI(n10127), .I0(state_timeout_counter[26]), 
            .I1(VCC_net), .CO(n10128));
    SB_CARRY sub_31_add_2_13 (.CI(n10112), .I0(state_timeout_counter[11]), 
            .I1(VCC_net), .CO(n10113));
    SB_LUT4 sub_31_add_2_12_lut (.I0(n1774), .I1(state_timeout_counter[10]), 
            .I2(VCC_net), .I3(n10111), .O(n12048)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_27_lut (.I0(GND_net), .I1(state_timeout_counter[25]), 
            .I2(VCC_net), .I3(n10126), .O(n506[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_12 (.CI(n10111), .I0(state_timeout_counter[10]), 
            .I1(VCC_net), .CO(n10112));
    SB_LUT4 sub_31_add_2_11_lut (.I0(n1774), .I1(state_timeout_counter[9]), 
            .I2(VCC_net), .I3(n10110), .O(n12049)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_27 (.CI(n10126), .I0(state_timeout_counter[25]), 
            .I1(VCC_net), .CO(n10127));
    SB_CARRY sub_31_add_2_11 (.CI(n10110), .I0(state_timeout_counter[9]), 
            .I1(VCC_net), .CO(n10111));
    SB_LUT4 sub_31_add_2_10_lut (.I0(GND_net), .I1(state_timeout_counter[8]), 
            .I2(VCC_net), .I3(n10109), .O(n506[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_26_lut (.I0(n1774), .I1(state_timeout_counter[24]), 
            .I2(VCC_net), .I3(n10125), .O(n12039)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_26 (.CI(n10125), .I0(state_timeout_counter[24]), 
            .I1(VCC_net), .CO(n10126));
    SB_LUT4 sub_31_add_2_25_lut (.I0(n1774), .I1(state_timeout_counter[23]), 
            .I2(VCC_net), .I3(n10124), .O(n12040)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_25 (.CI(n10124), .I0(state_timeout_counter[23]), 
            .I1(VCC_net), .CO(n10125));
    SB_LUT4 sub_31_add_2_24_lut (.I0(n1774), .I1(state_timeout_counter[22]), 
            .I2(VCC_net), .I3(n10123), .O(n12041)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_10 (.CI(n10109), .I0(state_timeout_counter[8]), 
            .I1(VCC_net), .CO(n10110));
    SB_LUT4 sub_31_add_2_9_lut (.I0(GND_net), .I1(state_timeout_counter[7]), 
            .I2(VCC_net), .I3(n10108), .O(n506[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_24 (.CI(n10123), .I0(state_timeout_counter[22]), 
            .I1(VCC_net), .CO(n10124));
    SB_DFFESR state_timeout_counter_i0_i8 (.Q(state_timeout_counter[8]), .C(SLM_CLK_c), 
            .E(n4491), .D(n506[8]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFF invert_55_i3 (.Q(INVERT_c_3), .C(SLM_CLK_c), .D(n968[3]));   // src/timing_controller.v(62[5] 131[12])
    SB_CARRY sub_31_add_2_9 (.CI(n10108), .I0(state_timeout_counter[7]), 
            .I1(VCC_net), .CO(n10109));
    SB_LUT4 sub_31_add_2_8_lut (.I0(GND_net), .I1(state_timeout_counter[6]), 
            .I2(VCC_net), .I3(n10107), .O(n506[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_23_lut (.I0(GND_net), .I1(state_timeout_counter[21]), 
            .I2(VCC_net), .I3(n10122), .O(n506[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_8 (.CI(n10107), .I0(state_timeout_counter[6]), 
            .I1(VCC_net), .CO(n10108));
    SB_DFFESR state_timeout_counter_i0_i7 (.Q(state_timeout_counter[7]), .C(SLM_CLK_c), 
            .E(n4491), .D(n506[7]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i6 (.Q(state_timeout_counter[6]), .C(SLM_CLK_c), 
            .E(n4491), .D(n506[6]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1880[2]), .R(n4806));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1880[1]), .R(n4806));   // src/timing_controller.v(56[8] 132[4])
    SB_CARRY sub_31_add_2_23 (.CI(n10122), .I0(state_timeout_counter[21]), 
            .I1(VCC_net), .CO(n10123));
    SB_LUT4 sub_31_add_2_7_lut (.I0(n10823), .I1(state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n10106), .O(n12054)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_DFF invert_55_i1 (.Q(buffer_switch_done), .C(SLM_CLK_c), .D(n13875));   // src/timing_controller.v(62[5] 131[12])
    SB_CARRY sub_31_add_2_7 (.CI(n10106), .I0(state_timeout_counter[5]), 
            .I1(VCC_net), .CO(n10107));
    SB_LUT4 sub_31_add_2_22_lut (.I0(n1774), .I1(state_timeout_counter[20]), 
            .I2(VCC_net), .I3(n10121), .O(n12042)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_6_lut (.I0(n1774), .I1(state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n10105), .O(n12106)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n4245));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6205_3_lut (.I0(state[0]), .I1(state[1]), .I2(state[2]), 
            .I3(GND_net), .O(n7568));
    defparam i6205_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_70 (.I0(n1774), .I1(n1879), .I2(GND_net), .I3(GND_net), 
            .O(n10823));   // src/timing_controller.v(62[5] 131[12])
    defparam i1_2_lut_adj_70.LUT_INIT = 16'h2222;
    SB_LUT4 i959_4_lut (.I0(state[3]), .I1(n2033), .I2(n7590), .I3(state[2]), 
            .O(n1951));   // src/timing_controller.v(56[8] 132[4])
    defparam i959_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i10384_2_lut (.I0(state[3]), .I1(n4192), .I2(GND_net), .I3(GND_net), 
            .O(n4491));   // src/timing_controller.v(62[5] 131[12])
    defparam i10384_2_lut.LUT_INIT = 16'h7777;
    SB_DFFE state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[0]));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFE state_i2 (.Q(state[2]), .C(SLM_CLK_c), .E(n4496), .D(state_3__N_80[2]));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFE state_i1 (.Q(state[1]), .C(SLM_CLK_c), .E(n4496), .D(state_3__N_80[1]));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFE state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[3]));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFE state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[4]));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFE state_timeout_counter_i0_i5 (.Q(state_timeout_counter[5]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[5]));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFE state_timeout_counter_i0_i9 (.Q(state_timeout_counter[9]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[9]));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFE state_timeout_counter_i0_i10 (.Q(state_timeout_counter[10]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[10]));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFE state_timeout_counter_i0_i12 (.Q(state_timeout_counter[12]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[12]));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFE state_timeout_counter_i0_i14 (.Q(state_timeout_counter[14]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[14]));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFE state_timeout_counter_i0_i15 (.Q(state_timeout_counter[15]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[15]));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFE state_timeout_counter_i0_i18 (.Q(state_timeout_counter[18]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[18]));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFE state_timeout_counter_i0_i19 (.Q(state_timeout_counter[19]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[19]));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFE state_timeout_counter_i0_i20 (.Q(state_timeout_counter[20]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[20]));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFE state_timeout_counter_i0_i22 (.Q(state_timeout_counter[22]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[22]));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFE state_timeout_counter_i0_i23 (.Q(state_timeout_counter[23]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[23]));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFE state_timeout_counter_i0_i24 (.Q(state_timeout_counter[24]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[24]));   // src/timing_controller.v(56[8] 132[4])
    SB_LUT4 i1_2_lut_3_lut (.I0(state[2]), .I1(state[0]), .I2(n63), .I3(GND_net), 
            .O(n10837));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i948_2_lut_3_lut (.I0(state[0]), .I1(n63), .I2(state[1]), 
            .I3(GND_net), .O(n2033));   // src/timing_controller.v(56[8] 132[4])
    defparam i948_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 mux_343_Mux_3_i15_4_lut_4_lut (.I0(state[2]), .I1(state[0]), 
            .I2(state[1]), .I3(state[3]), .O(n968[3]));
    defparam mux_343_Mux_3_i15_4_lut_4_lut.LUT_INIT = 16'h01a0;
    SB_LUT4 i6_2_lut (.I0(state_timeout_counter[9]), .I1(state_timeout_counter[12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // src/timing_controller.v(84[17:45])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut (.I0(state_timeout_counter[17]), .I1(state_timeout_counter[1]), 
            .I2(state_timeout_counter[24]), .I3(state_timeout_counter[4]), 
            .O(n52));   // src/timing_controller.v(84[17:45])
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(state_timeout_counter[29]), .I1(state_timeout_counter[3]), 
            .I2(state_timeout_counter[13]), .I3(state_timeout_counter[31]), 
            .O(n56));   // src/timing_controller.v(84[17:45])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(state_timeout_counter[19]), .I1(state_timeout_counter[5]), 
            .I2(state_timeout_counter[22]), .I3(state_timeout_counter[6]), 
            .O(n54));   // src/timing_controller.v(84[17:45])
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(state_timeout_counter[10]), .I1(state_timeout_counter[15]), 
            .I2(state_timeout_counter[20]), .I3(state_timeout_counter[23]), 
            .O(n55));   // src/timing_controller.v(84[17:45])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(state_timeout_counter[27]), .I1(state_timeout_counter[7]), 
            .I2(state_timeout_counter[30]), .I3(state_timeout_counter[14]), 
            .O(n53));   // src/timing_controller.v(84[17:45])
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(state_timeout_counter[8]), .I1(state_timeout_counter[11]), 
            .I2(state_timeout_counter[16]), .I3(state_timeout_counter[21]), 
            .O(n50));   // src/timing_controller.v(84[17:45])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(state_timeout_counter[25]), .I1(n52), .I2(n38), 
            .I3(state_timeout_counter[26]), .O(n58));   // src/timing_controller.v(84[17:45])
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30_4_lut (.I0(n53), .I1(n55), .I2(n54), .I3(n56), .O(n62));   // src/timing_controller.v(84[17:45])
    defparam i30_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(state_timeout_counter[0]), .I1(state_timeout_counter[18]), 
            .I2(state_timeout_counter[28]), .I3(state_timeout_counter[2]), 
            .O(n49));   // src/timing_controller.v(84[17:45])
    defparam i17_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i31_4_lut (.I0(n49), .I1(n62), .I2(n58), .I3(n50), .O(n63));   // src/timing_controller.v(84[17:45])
    defparam i31_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_71 (.I0(state[3]), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n10831));
    defparam i1_2_lut_adj_71.LUT_INIT = 16'hbbbb;
    SB_LUT4 i6207_3_lut (.I0(n63), .I1(state[1]), .I2(state[2]), .I3(GND_net), 
            .O(n7570));
    defparam i6207_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 state_3__I_0_59_Mux_0_i7_4_lut (.I0(state[1]), .I1(n63), .I2(state[2]), 
            .I3(state[0]), .O(n7));   // src/timing_controller.v(62[5] 131[12])
    defparam state_3__I_0_59_Mux_0_i7_4_lut.LUT_INIT = 16'hc535;
    SB_LUT4 state_3__I_0_59_Mux_0_i15_4_lut (.I0(n7), .I1(n7570), .I2(state[3]), 
            .I3(state[0]), .O(state_3__N_80[0]));   // src/timing_controller.v(62[5] 131[12])
    defparam state_3__I_0_59_Mux_0_i15_4_lut.LUT_INIT = 16'hfa3a;
    SB_DFFESR invert_55_i2 (.Q(UPDATE_c_2), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n12202), .R(n5));   // src/timing_controller.v(62[5] 131[12])
    SB_LUT4 i1_2_lut_3_lut_adj_72 (.I0(n7568), .I1(state[3]), .I2(n63), 
            .I3(GND_net), .O(n4496));
    defparam i1_2_lut_3_lut_adj_72.LUT_INIT = 16'hdfdf;
    SB_LUT4 mux_898_i1_4_lut (.I0(n1880[0]), .I1(state[1]), .I2(n1951), 
            .I3(n10814), .O(n1952[0]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_898_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 mux_890_i1_3_lut (.I0(n12036), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[0]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i1_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10438_2_lut (.I0(state[3]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // src/timing_controller.v(56[8] 132[4])
    defparam i10438_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[3]), .I1(n63), .I2(state[1]), .I3(state[2]), 
            .O(n10833));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(state[0]), .I1(n63), .I2(state[3]), 
            .I3(state[2]), .O(n10814));   // src/timing_controller.v(56[8] 132[4])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 state_3__I_0_59_Mux_2_i15_4_lut (.I0(state[1]), .I1(state[2]), 
            .I2(state[3]), .I3(state[0]), .O(state_3__N_80[2]));   // src/timing_controller.v(62[5] 131[12])
    defparam state_3__I_0_59_Mux_2_i15_4_lut.LUT_INIT = 16'hc2ce;
    SB_LUT4 i10442_3_lut_4_lut (.I0(state[3]), .I1(n4192), .I2(n1951), 
            .I3(n10823), .O(n4809));
    defparam i10442_3_lut_4_lut.LUT_INIT = 16'h7077;
    SB_LUT4 state_3__I_0_59_Mux_1_i15_4_lut_4_lut (.I0(state[0]), .I1(state[1]), 
            .I2(state[3]), .I3(n10837), .O(state_3__N_80[1]));   // src/timing_controller.v(62[5] 131[12])
    defparam state_3__I_0_59_Mux_1_i15_4_lut_4_lut.LUT_INIT = 16'hc6f6;
    SB_LUT4 i1_2_lut_3_lut_adj_73 (.I0(state[2]), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n4192));
    defparam i1_2_lut_3_lut_adj_73.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_890_i4_3_lut (.I0(n12050), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[3]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9121_4_lut (.I0(n12106), .I1(state[1]), .I2(n1879), .I3(n1951), 
            .O(n1952[4]));   // src/timing_controller.v(62[5] 131[12])
    defparam i9121_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_898_i6_3_lut (.I0(n12054), .I1(state[1]), .I2(n1951), 
            .I3(GND_net), .O(n1952[5]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_898_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_890_i10_3_lut (.I0(n12049), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[9]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i10_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i11_3_lut (.I0(n12048), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[10]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i11_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i13_3_lut (.I0(n12047), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[12]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i13_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i15_3_lut (.I0(n12046), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[14]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i15_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i16_3_lut (.I0(n12045), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[15]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i16_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i19_3_lut (.I0(n12044), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[18]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i19_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i20_3_lut (.I0(n12043), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[19]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i21_3_lut (.I0(n12042), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[20]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i21_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i23_3_lut (.I0(n12041), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[22]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i23_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i24_3_lut (.I0(n12040), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[23]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i3423_2_lut_3_lut (.I0(state[3]), .I1(n4192), .I2(n1951), 
            .I3(GND_net), .O(n4806));   // src/timing_controller.v(56[8] 132[4])
    defparam i3423_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 mux_890_i25_3_lut (.I0(n12039), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[24]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i25_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10364_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n12202));   // src/timing_controller.v(62[5] 131[12])
    defparam i10364_2_lut.LUT_INIT = 16'h9999;
    
endmodule
//
// Verilog Description of module bluejay_data
//

module bluejay_data (dc32_fifo_almost_full, n771, dc32_fifo_almost_empty, 
            bluejay_data_out_31__N_736, buffer_switch_done_latched, GND_net, 
            DEBUG_9_c, SLM_CLK_c, DATA19_c, buffer_switch_done, n4937, 
            DATA18_c, n4936, DATA17_c, n6112, DEBUG_6_c, DATA15_c, 
            DATA14_c, DATA13_c, DATA12_c, n843, VCC_net, DATA11_c, 
            DATA10_c, SYNC_c, bluejay_data_out_31__N_737, n10277, DATA9_c, 
            DATA8_c, DATA7_c, DATA6_c, \rd_sig_diff0_w[1] , get_next_word, 
            \rd_sig_diff0_w[0] , \rd_sig_diff0_w[2] , n10873, n10877, 
            \aempty_flag_impl.ae_flag_nxt_w , DATA5_c, DATA20_c, \fifo_data_out[4] , 
            \fifo_data_out[5] , \fifo_data_out[6] , \fifo_data_out[7] , 
            \fifo_data_out[11] , \fifo_data_out[10] , \fifo_data_out[3] , 
            \fifo_data_out[15] , \fifo_data_out[14] , \fifo_data_out[13] , 
            \fifo_data_out[12] , \fifo_data_out[9] , \fifo_data_out[8] ) /* synthesis syn_module_defined=1 */ ;
    input dc32_fifo_almost_full;
    output n771;
    input dc32_fifo_almost_empty;
    output bluejay_data_out_31__N_736;
    input buffer_switch_done_latched;
    input GND_net;
    output DEBUG_9_c;
    input SLM_CLK_c;
    output DATA19_c;
    input buffer_switch_done;
    input n4937;
    output DATA18_c;
    input n4936;
    output DATA17_c;
    input n6112;
    output DEBUG_6_c;
    output DATA15_c;
    output DATA14_c;
    output DATA13_c;
    output DATA12_c;
    output n843;
    input VCC_net;
    output DATA11_c;
    output DATA10_c;
    output SYNC_c;
    output bluejay_data_out_31__N_737;
    input n10277;
    output DATA9_c;
    output DATA8_c;
    output DATA7_c;
    output DATA6_c;
    input \rd_sig_diff0_w[1] ;
    output get_next_word;
    input \rd_sig_diff0_w[0] ;
    input \rd_sig_diff0_w[2] ;
    input n10873;
    input n10877;
    output \aempty_flag_impl.ae_flag_nxt_w ;
    output DATA5_c;
    output DATA20_c;
    input \fifo_data_out[4] ;
    input \fifo_data_out[5] ;
    input \fifo_data_out[6] ;
    input \fifo_data_out[7] ;
    input \fifo_data_out[11] ;
    input \fifo_data_out[10] ;
    input \fifo_data_out[3] ;
    input \fifo_data_out[15] ;
    input \fifo_data_out[14] ;
    input \fifo_data_out[13] ;
    input \fifo_data_out[12] ;
    input \fifo_data_out[9] ;
    input \fifo_data_out[8] ;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [15:0]n828;
    
    wire n891, bluejay_data_out_31__N_735, n3033, n895, valid_N_740, 
        n6575, n1, n4, n4370, n4704, n4938;
    wire [10:0]v_counter_10__N_715;
    
    wire n4408;
    wire [10:0]v_counter;   // src/bluejay_data.v(51[12:21])
    
    wire n6071, n6041, n6023, n6022, n10969, n10967, n4_adj_46, 
        n20, n10989;
    wire [7:0]state_timeout_counter;   // src/bluejay_data.v(52[11:32])
    
    wire n10891, n13, n10977, n1291, n27, n10594, n4228, n10154, 
        n10153, n10152, n10151, n12, n10306, n10307, n10240, n10150, 
        n10149, n3031, n10148, n10147, n5886, n10146, n5869, n10145;
    wire [8:0]n62;
    
    wire n10089, n10088, n1_adj_47, n10085, n1_adj_48, n10083, n10084, 
        n10086, n10087, bluejay_data_out_31__N_734, n3035, n3029, 
        n1_adj_49, n5557, n1_adj_50, n1_adj_51, n5475, n5308, n12_adj_52, 
        n5291, n15, n5258, n4679, n4710, n10708, n4876, n7469, 
        n5058;
    
    SB_LUT4 reduce_or_325_i1_4_lut (.I0(dc32_fifo_almost_full), .I1(n771), 
            .I2(n828[5]), .I3(n828[4]), .O(n891));   // src/bluejay_data.v(66[9] 121[16])
    defparam reduce_or_325_i1_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 i1_4_lut (.I0(dc32_fifo_almost_empty), .I1(bluejay_data_out_31__N_735), 
            .I2(bluejay_data_out_31__N_736), .I3(buffer_switch_done_latched), 
            .O(n3033));   // src/bluejay_data.v(43[15:31])
    defparam i1_4_lut.LUT_INIT = 16'hccdc;
    SB_LUT4 i1_2_lut (.I0(bluejay_data_out_31__N_736), .I1(dc32_fifo_almost_empty), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_DFFN valid_56 (.Q(DEBUG_9_c), .C(SLM_CLK_c), .D(valid_N_740));   // src/bluejay_data.v(126[8] 148[4])
    SB_LUT4 i1_2_lut_3_lut (.I0(buffer_switch_done_latched), .I1(n6575), 
            .I2(n1), .I3(GND_net), .O(n4));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3321_3_lut_4_lut (.I0(buffer_switch_done_latched), .I1(n6575), 
            .I2(bluejay_data_out_31__N_735), .I3(n4370), .O(n4704));   // src/bluejay_data.v(66[9] 121[16])
    defparam i3321_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_DFFN bluejay_data_out_i4 (.Q(DATA19_c), .C(SLM_CLK_c), .D(n4938));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFESR v_counter_i1 (.Q(v_counter[1]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[1]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i2 (.Q(v_counter[2]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[2]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i3 (.Q(v_counter[3]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[3]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFN bluejay_data_out_i3 (.Q(DATA18_c), .C(SLM_CLK_c), .D(n4937));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFESR v_counter_i4 (.Q(v_counter[4]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[4]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i5 (.Q(v_counter[5]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[5]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i6 (.Q(v_counter[6]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[6]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i7 (.Q(v_counter[7]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[7]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESS v_counter_i8 (.Q(v_counter[8]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[8]), .S(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i9 (.Q(v_counter[9]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[9]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESS v_counter_i10 (.Q(v_counter[10]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[10]), .S(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFN bluejay_data_out_i2 (.Q(DATA17_c), .C(SLM_CLK_c), .D(n4936));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i1 (.Q(DEBUG_6_c), .C(SLM_CLK_c), .D(n6112));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i16 (.Q(DATA15_c), .C(SLM_CLK_c), .D(n6071));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i15 (.Q(DATA14_c), .C(SLM_CLK_c), .D(n6041));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i14 (.Q(DATA13_c), .C(SLM_CLK_c), .D(n6023));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i13 (.Q(DATA12_c), .C(SLM_CLK_c), .D(n6022));   // src/bluejay_data.v(126[8] 148[4])
    SB_LUT4 i9132_4_lut (.I0(v_counter[8]), .I1(v_counter[4]), .I2(v_counter[5]), 
            .I3(v_counter[3]), .O(n10969));
    defparam i9132_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9130_4_lut (.I0(v_counter[2]), .I1(v_counter[6]), .I2(v_counter[7]), 
            .I3(v_counter[9]), .O(n10967));
    defparam i9130_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_43 (.I0(dc32_fifo_almost_full), .I1(n843), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_46));
    defparam i1_2_lut_adj_43.LUT_INIT = 16'h4444;
    SB_LUT4 i9151_4_lut (.I0(n10967), .I1(n20), .I2(n10969), .I3(v_counter[10]), 
            .O(n10989));
    defparam i9151_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9055_2_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[5]), 
            .I2(GND_net), .I3(GND_net), .O(n10891));
    defparam i9055_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9139_4_lut (.I0(state_timeout_counter[3]), .I1(state_timeout_counter[2]), 
            .I2(state_timeout_counter[4]), .I3(n13), .O(n10977));
    defparam i9139_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(n828[9]), .I1(n828[4]), .I2(n843), .I3(GND_net), 
            .O(n1291));   // src/bluejay_data.v(66[9] 121[16])
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_44 (.I0(state_timeout_counter[0]), .I1(n10989), 
            .I2(n4_adj_46), .I3(n828[9]), .O(n27));
    defparam i1_4_lut_adj_44.LUT_INIT = 16'ha2a0;
    SB_LUT4 i1_4_lut_adj_45 (.I0(n828[2]), .I1(n27), .I2(n10977), .I3(n10891), 
            .O(n10594));
    defparam i1_4_lut_adj_45.LUT_INIT = 16'haaae;
    SB_LUT4 i1_3_lut (.I0(dc32_fifo_almost_full), .I1(n843), .I2(n771), 
            .I3(GND_net), .O(n4228));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 sub_118_add_2_12_lut (.I0(GND_net), .I1(v_counter[10]), .I2(VCC_net), 
            .I3(n10154), .O(v_counter_10__N_715[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_118_add_2_11_lut (.I0(GND_net), .I1(v_counter[9]), .I2(VCC_net), 
            .I3(n10153), .O(v_counter_10__N_715[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_11 (.CI(n10153), .I0(v_counter[9]), .I1(VCC_net), 
            .CO(n10154));
    SB_LUT4 sub_118_add_2_10_lut (.I0(GND_net), .I1(v_counter[8]), .I2(VCC_net), 
            .I3(n10152), .O(v_counter_10__N_715[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 equal_1263_i20_2_lut (.I0(v_counter[0]), .I1(v_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n20));   // src/bluejay_data.v(106[21:49])
    defparam equal_1263_i20_2_lut.LUT_INIT = 16'hdddd;
    SB_CARRY sub_118_add_2_10 (.CI(n10152), .I0(v_counter[8]), .I1(VCC_net), 
            .CO(n10153));
    SB_LUT4 sub_118_add_2_9_lut (.I0(GND_net), .I1(v_counter[7]), .I2(VCC_net), 
            .I3(n10151), .O(v_counter_10__N_715[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_4_lut (.I0(v_counter[8]), .I1(v_counter[7]), .I2(v_counter[4]), 
            .I3(v_counter[3]), .O(n12));   // src/bluejay_data.v(108[25:41])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY sub_118_add_2_9 (.CI(n10151), .I0(v_counter[7]), .I1(VCC_net), 
            .CO(n10152));
    SB_LUT4 i6_4_lut (.I0(v_counter[5]), .I1(n12), .I2(v_counter[2]), 
            .I3(v_counter[6]), .O(n10306));   // src/bluejay_data.v(108[25:41])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n828[9]), .I1(n10306), .I2(n771), .I3(n10307), 
            .O(n10240));   // src/bluejay_data.v(66[9] 121[16])
    defparam i2_4_lut.LUT_INIT = 16'h0a08;
    SB_LUT4 sub_118_add_2_8_lut (.I0(GND_net), .I1(v_counter[6]), .I2(VCC_net), 
            .I3(n10150), .O(v_counter_10__N_715[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_8 (.CI(n10150), .I0(v_counter[6]), .I1(VCC_net), 
            .CO(n10151));
    SB_LUT4 sub_118_add_2_7_lut (.I0(GND_net), .I1(v_counter[5]), .I2(VCC_net), 
            .I3(n10149), .O(v_counter_10__N_715[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_7 (.CI(n10149), .I0(v_counter[5]), .I1(VCC_net), 
            .CO(n10150));
    SB_LUT4 i1664_4_lut (.I0(buffer_switch_done_latched), .I1(n10240), .I2(n828[5]), 
            .I3(dc32_fifo_almost_full), .O(n3031));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1664_4_lut.LUT_INIT = 16'hccdc;
    SB_LUT4 sub_118_add_2_6_lut (.I0(GND_net), .I1(v_counter[4]), .I2(VCC_net), 
            .I3(n10148), .O(v_counter_10__N_715[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_6 (.CI(n10148), .I0(v_counter[4]), .I1(VCC_net), 
            .CO(n10149));
    SB_LUT4 sub_118_add_2_5_lut (.I0(GND_net), .I1(v_counter[3]), .I2(VCC_net), 
            .I3(n10147), .O(v_counter_10__N_715[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFN bluejay_data_out_i12 (.Q(DATA11_c), .C(SLM_CLK_c), .D(n5886));   // src/bluejay_data.v(126[8] 148[4])
    SB_CARRY sub_118_add_2_5 (.CI(n10147), .I0(v_counter[3]), .I1(VCC_net), 
            .CO(n10148));
    SB_LUT4 sub_118_add_2_4_lut (.I0(GND_net), .I1(v_counter[2]), .I2(VCC_net), 
            .I3(n10146), .O(v_counter_10__N_715[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_4 (.CI(n10146), .I0(v_counter[2]), .I1(VCC_net), 
            .CO(n10147));
    SB_DFFN bluejay_data_out_i11 (.Q(DATA10_c), .C(SLM_CLK_c), .D(n5869));   // src/bluejay_data.v(126[8] 148[4])
    SB_LUT4 sub_118_add_2_3_lut (.I0(GND_net), .I1(v_counter[1]), .I2(VCC_net), 
            .I3(n10145), .O(v_counter_10__N_715[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_3 (.CI(n10145), .I0(v_counter[1]), .I1(VCC_net), 
            .CO(n10146));
    SB_LUT4 sub_118_add_2_2_lut (.I0(GND_net), .I1(v_counter[0]), .I2(n771), 
            .I3(VCC_net), .O(v_counter_10__N_715[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_2 (.CI(VCC_net), .I0(v_counter[0]), .I1(n771), 
            .CO(n10145));
    SB_LUT4 sub_116_add_2_9_lut (.I0(GND_net), .I1(state_timeout_counter[7]), 
            .I2(VCC_net), .I3(n10089), .O(n62[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_46 (.I0(n828[9]), .I1(buffer_switch_done), .I2(GND_net), 
            .I3(GND_net), .O(n4408));
    defparam i1_2_lut_adj_46.LUT_INIT = 16'heeee;
    SB_LUT4 sub_116_add_2_8_lut (.I0(GND_net), .I1(state_timeout_counter[6]), 
            .I2(VCC_net), .I3(n10088), .O(n62[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_116_add_2_8 (.CI(n10088), .I0(state_timeout_counter[6]), 
            .I1(VCC_net), .CO(n10089));
    SB_LUT4 sub_116_add_2_5_lut (.I0(n1291), .I1(state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n10085), .O(n1_adj_47)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_116_add_2_3_lut (.I0(n1291), .I1(state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n10083), .O(n1_adj_48)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_116_add_2_3 (.CI(n10083), .I0(state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n10084));
    SB_CARRY sub_116_add_2_6 (.CI(n10086), .I0(state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n10087));
    SB_DFFN sync_58 (.Q(SYNC_c), .C(SLM_CLK_c), .D(bluejay_data_out_31__N_734));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFSR state_FSM_i10 (.Q(n828[9]), .C(SLM_CLK_c), .D(n3035), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i9 (.Q(bluejay_data_out_31__N_737), .C(SLM_CLK_c), 
            .D(n895), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i8 (.Q(bluejay_data_out_31__N_736), .C(SLM_CLK_c), 
            .D(n3033), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i7 (.Q(bluejay_data_out_31__N_735), .C(SLM_CLK_c), 
            .D(n891), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i6 (.Q(n828[5]), .C(SLM_CLK_c), .D(n3031), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i5 (.Q(n828[4]), .C(SLM_CLK_c), .D(n3029), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i4 (.Q(bluejay_data_out_31__N_734), .C(SLM_CLK_c), 
            .D(n4228), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i3 (.Q(n828[2]), .C(SLM_CLK_c), .D(n10594), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i2 (.Q(n843), .C(SLM_CLK_c), .D(n10277), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_CARRY sub_116_add_2_5 (.CI(n10085), .I0(state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n10086));
    SB_LUT4 sub_116_add_2_7_lut (.I0(n1291), .I1(state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n10087), .O(n1_adj_49)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_DFFN bluejay_data_out_i10 (.Q(DATA9_c), .C(SLM_CLK_c), .D(n5557));   // src/bluejay_data.v(126[8] 148[4])
    SB_CARRY sub_116_add_2_7 (.CI(n10087), .I0(state_timeout_counter[5]), 
            .I1(VCC_net), .CO(n10088));
    SB_LUT4 sub_116_add_2_6_lut (.I0(n1291), .I1(state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n10086), .O(n1_adj_50)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_116_add_2_2_lut (.I0(n1291), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n1_adj_51)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_116_add_2_4_lut (.I0(n1291), .I1(state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n10084), .O(n1)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_116_add_2_2 (.CI(VCC_net), .I0(state_timeout_counter[0]), 
            .I1(GND_net), .CO(n10083));
    SB_CARRY sub_116_add_2_4 (.CI(n10084), .I0(state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n10085));
    SB_DFFN bluejay_data_out_i9 (.Q(DATA8_c), .C(SLM_CLK_c), .D(n5475));   // src/bluejay_data.v(126[8] 148[4])
    SB_LUT4 equal_117_i13_2_lut (.I0(state_timeout_counter[6]), .I1(state_timeout_counter[7]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // src/bluejay_data.v(106[21:49])
    defparam equal_117_i13_2_lut.LUT_INIT = 16'heeee;
    SB_DFFN bluejay_data_out_i8 (.Q(DATA7_c), .C(SLM_CLK_c), .D(n5308));   // src/bluejay_data.v(126[8] 148[4])
    SB_LUT4 i5_4_lut_adj_47 (.I0(state_timeout_counter[3]), .I1(n13), .I2(state_timeout_counter[1]), 
            .I3(state_timeout_counter[2]), .O(n12_adj_52));   // src/bluejay_data.v(106[21:49])
    defparam i5_4_lut_adj_47.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_48 (.I0(state_timeout_counter[4]), .I1(n12_adj_52), 
            .I2(state_timeout_counter[5]), .I3(state_timeout_counter[0]), 
            .O(n771));   // src/bluejay_data.v(106[21:49])
    defparam i6_4_lut_adj_48.LUT_INIT = 16'hfeff;
    SB_DFFN bluejay_data_out_i7 (.Q(DATA6_c), .C(SLM_CLK_c), .D(n5291));   // src/bluejay_data.v(126[8] 148[4])
    SB_LUT4 i1_3_lut_adj_49 (.I0(\rd_sig_diff0_w[1] ), .I1(get_next_word), 
            .I2(\rd_sig_diff0_w[0] ), .I3(GND_net), .O(n15));   // src/fifo_dc_32_lut_gen.v(233[30:44])
    defparam i1_3_lut_adj_49.LUT_INIT = 16'h5d5d;
    SB_LUT4 i5_4_lut_adj_50 (.I0(\rd_sig_diff0_w[2] ), .I1(n10873), .I2(n15), 
            .I3(n10877), .O(\aempty_flag_impl.ae_flag_nxt_w ));   // src/fifo_dc_32_lut_gen.v(233[30:44])
    defparam i5_4_lut_adj_50.LUT_INIT = 16'h0010;
    SB_DFFN bluejay_data_out_i6 (.Q(DATA5_c), .C(SLM_CLK_c), .D(n5258));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFESS state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(SLM_CLK_c), 
            .E(n4370), .D(n1_adj_48), .S(n4679));   // src/bluejay_data.v(56[8] 123[4])
    SB_LUT4 i1_3_lut_4_lut (.I0(buffer_switch_done_latched), .I1(n771), 
            .I2(n828[9]), .I3(bluejay_data_out_31__N_737), .O(n3035));   // src/bluejay_data.v(62[9] 65[12])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hff40;
    SB_DFFESS state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(SLM_CLK_c), 
            .E(n4370), .D(n4), .S(n4710));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESS state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(SLM_CLK_c), 
            .E(n4370), .D(n1_adj_47), .S(n4704));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESS state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(SLM_CLK_c), 
            .E(n4370), .D(n1_adj_50), .S(n10708));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFN get_next_word_57 (.Q(get_next_word), .C(SLM_CLK_c), .D(n4876));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFESS state_timeout_counter_i0_i5 (.Q(state_timeout_counter[5]), .C(SLM_CLK_c), 
            .E(n4370), .D(n1_adj_49), .S(n4704));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR state_timeout_counter_i0_i6 (.Q(state_timeout_counter[6]), .C(SLM_CLK_c), 
            .E(n4370), .D(n62[6]), .R(n7469));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR state_timeout_counter_i0_i7 (.Q(state_timeout_counter[7]), .C(SLM_CLK_c), 
            .E(n4370), .D(n62[7]), .R(n7469));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESS state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(SLM_CLK_c), 
            .E(n4370), .D(n1_adj_51), .S(n4679));   // src/bluejay_data.v(56[8] 123[4])
    SB_LUT4 i1662_3_lut_4_lut (.I0(buffer_switch_done_latched), .I1(n771), 
            .I2(bluejay_data_out_31__N_734), .I3(n828[4]), .O(n3029));   // src/bluejay_data.v(62[9] 65[12])
    defparam i1662_3_lut_4_lut.LUT_INIT = 16'hf4f0;
    SB_LUT4 i1_2_lut_adj_51 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_737), 
            .I2(GND_net), .I3(GND_net), .O(valid_N_740));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1_2_lut_adj_51.LUT_INIT = 16'heeee;
    SB_DFFN bluejay_data_out_i5 (.Q(DATA20_c), .C(SLM_CLK_c), .D(n5058));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFESR v_counter_i0 (.Q(v_counter[0]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[0]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_LUT4 i10434_3_lut (.I0(buffer_switch_done_latched), .I1(buffer_switch_done), 
            .I2(n6575), .I3(GND_net), .O(n4370));   // src/bluejay_data.v(61[10] 122[8])
    defparam i10434_3_lut.LUT_INIT = 16'h2323;
    SB_LUT4 i3296_2_lut (.I0(n4370), .I1(bluejay_data_out_31__N_734), .I2(GND_net), 
            .I3(GND_net), .O(n4679));   // src/bluejay_data.v(56[8] 123[4])
    defparam i3296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_52 (.I0(n828[2]), .I1(n828[5]), .I2(bluejay_data_out_31__N_736), 
            .I3(GND_net), .O(n6575));   // src/bluejay_data.v(66[9] 121[16])
    defparam i2_3_lut_adj_52.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_53 (.I0(n4370), .I1(bluejay_data_out_31__N_737), 
            .I2(GND_net), .I3(GND_net), .O(n4710));   // src/bluejay_data.v(61[10] 122[8])
    defparam i1_2_lut_adj_53.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_54 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_737), 
            .I2(\fifo_data_out[4] ), .I3(GND_net), .O(n5058));
    defparam i1_2_lut_3_lut_adj_54.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_55 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_737), 
            .I2(\fifo_data_out[5] ), .I3(GND_net), .O(n5258));
    defparam i1_2_lut_3_lut_adj_55.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_56 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_737), 
            .I2(\fifo_data_out[6] ), .I3(GND_net), .O(n5291));
    defparam i1_2_lut_3_lut_adj_56.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_57 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_737), 
            .I2(\fifo_data_out[7] ), .I3(GND_net), .O(n5308));
    defparam i1_2_lut_3_lut_adj_57.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_58 (.I0(buffer_switch_done_latched), .I1(buffer_switch_done), 
            .I2(GND_net), .I3(GND_net), .O(n10708));   // src/bluejay_data.v(61[10] 122[8])
    defparam i1_2_lut_adj_58.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_59 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_735), 
            .I2(GND_net), .I3(GND_net), .O(n4876));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1_2_lut_adj_59.LUT_INIT = 16'heeee;
    SB_LUT4 i10405_2_lut (.I0(n4370), .I1(n1291), .I2(GND_net), .I3(GND_net), 
            .O(n7469));
    defparam i10405_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_60 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_737), 
            .I2(\fifo_data_out[11] ), .I3(GND_net), .O(n5886));
    defparam i1_2_lut_3_lut_adj_60.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_61 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_737), 
            .I2(\fifo_data_out[10] ), .I3(GND_net), .O(n5869));
    defparam i1_2_lut_3_lut_adj_61.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_62 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_737), 
            .I2(\fifo_data_out[3] ), .I3(GND_net), .O(n4938));
    defparam i1_2_lut_3_lut_adj_62.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_3_lut_4_lut_adj_63 (.I0(v_counter[9]), .I1(v_counter[0]), 
            .I2(v_counter[1]), .I3(v_counter[10]), .O(n10307));   // src/bluejay_data.v(108[25:41])
    defparam i1_3_lut_4_lut_adj_63.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut_adj_64 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_737), 
            .I2(\fifo_data_out[15] ), .I3(GND_net), .O(n6071));
    defparam i1_2_lut_3_lut_adj_64.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_65 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_737), 
            .I2(\fifo_data_out[14] ), .I3(GND_net), .O(n6041));
    defparam i1_2_lut_3_lut_adj_65.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_66 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_737), 
            .I2(\fifo_data_out[13] ), .I3(GND_net), .O(n6023));
    defparam i1_2_lut_3_lut_adj_66.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_67 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_737), 
            .I2(\fifo_data_out[12] ), .I3(GND_net), .O(n6022));
    defparam i1_2_lut_3_lut_adj_67.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_68 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_737), 
            .I2(\fifo_data_out[9] ), .I3(GND_net), .O(n5557));
    defparam i1_2_lut_3_lut_adj_68.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_69 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_737), 
            .I2(\fifo_data_out[8] ), .I3(GND_net), .O(n5475));
    defparam i1_2_lut_3_lut_adj_69.LUT_INIT = 16'he0e0;
    
endmodule
//
// Verilog Description of module fifo_dc_32_lut_gen2
//

module fifo_dc_32_lut_gen2 (\rd_addr_r[0] , \REG.mem_14_5 , \REG.mem_15_5 , 
            \dc32_fifo_data_in[6] , dc32_fifo_almost_full, FIFO_CLK_c, 
            reset_per_frame, \REG.mem_13_5 , \REG.mem_12_5 , \dc32_fifo_data_in[5] , 
            \dc32_fifo_data_in[4] , \REG.mem_31_0 , GND_net, \dc32_fifo_data_in[3] , 
            \REG.mem_55_13 , \dc32_fifo_data_in[2] , \REG.mem_38_7 , \REG.mem_39_7 , 
            \REG.mem_36_7 , \REG.mem_37_7 , \REG.mem_16_8 , \REG.mem_18_8 , 
            \REG.mem_3_13 , \REG.mem_57_6 , \dc32_fifo_data_in[1] , \REG.mem_63_11 , 
            \dc32_fifo_data_in[0] , \REG.mem_35_0 , t_rd_fifo_en_w, \REG.out_raw[0] , 
            SLM_CLK_c, \REG.mem_55_10 , n62, n30, \REG.mem_31_3 , 
            \REG.mem_48_7 , \REG.mem_50_7 , \REG.mem_55_7 , \REG.mem_48_10 , 
            \REG.mem_50_10 , wr_grey_sync_r, \wr_addr_nxt_c[5] , \REG.mem_23_8 , 
            \REG.mem_25_5 , \rd_grey_sync_r[0] , \REG.mem_25_15 , \REG.mem_14_12 , 
            \REG.mem_15_12 , DEBUG_3_c, \REG.mem_13_12 , \REG.mem_12_12 , 
            \aempty_flag_impl.ae_flag_nxt_w , dc32_fifo_almost_empty, \REG.mem_6_1 , 
            \REG.mem_7_1 , \REG.mem_5_1 , \REG.mem_4_1 , \REG.mem_57_9 , 
            \REG.mem_35_3 , \REG.mem_46_1 , \REG.mem_47_1 , \REG.mem_45_1 , 
            \REG.mem_44_1 , \REG.mem_25_2 , \dc32_fifo_data_in[15] , \dc32_fifo_data_in[14] , 
            \dc32_fifo_data_in[13] , \REG.mem_3_11 , \REG.mem_31_2 , \REG.mem_50_12 , 
            \dc32_fifo_data_in[12] , \REG.mem_6_11 , \REG.mem_7_11 , \REG.mem_5_11 , 
            \REG.mem_4_11 , \dc32_fifo_data_in[11] , \REG.mem_48_12 , 
            \REG.mem_3_4 , \REG.mem_14_8 , \REG.mem_15_8 , \REG.mem_8_14 , 
            \REG.mem_9_14 , \dc32_fifo_data_in[10] , \REG.mem_10_14 , 
            \REG.mem_11_14 , \REG.mem_63_6 , \REG.mem_13_8 , \REG.mem_12_8 , 
            \REG.mem_14_14 , \REG.mem_15_14 , \dc32_fifo_data_in[9] , 
            \dc32_fifo_data_in[8] , \REG.mem_3_1 , \dc32_fifo_data_in[7] , 
            \REG.mem_12_14 , \REG.mem_13_14 , \REG.mem_42_8 , \REG.mem_43_8 , 
            \REG.mem_41_8 , \REG.mem_40_8 , \REG.mem_18_12 , \REG.mem_16_12 , 
            \REG.mem_31_15 , \REG.mem_38_3 , \REG.mem_39_3 , \REG.mem_37_3 , 
            \REG.mem_36_3 , \REG.mem_42_3 , \REG.mem_43_3 , \REG.mem_14_7 , 
            \REG.mem_15_7 , \REG.mem_13_7 , \REG.mem_12_7 , \REG.mem_41_3 , 
            \REG.mem_40_3 , \REG.mem_57_0 , \REG.mem_10_11 , \REG.mem_11_11 , 
            \REG.mem_9_11 , \REG.mem_8_11 , \REG.mem_63_12 , \REG.mem_55_12 , 
            \REG.mem_35_15 , \REG.mem_3_15 , \wr_addr_nxt_c[3] , \REG.mem_50_9 , 
            \REG.mem_48_9 , \REG.mem_46_8 , \REG.mem_47_8 , \REG.mem_46_3 , 
            \REG.mem_47_3 , \REG.mem_45_8 , \REG.mem_44_8 , \REG.mem_16_2 , 
            \REG.mem_10_9 , \REG.mem_11_9 , \REG.mem_45_3 , \REG.mem_44_3 , 
            \REG.mem_25_7 , \REG.mem_23_12 , \REG.mem_18_2 , \REG.mem_38_0 , 
            \REG.mem_39_0 , \REG.mem_31_13 , \REG.mem_37_0 , \REG.mem_36_0 , 
            \REG.mem_18_6 , \REG.mem_16_6 , \REG.mem_9_9 , \REG.mem_8_9 , 
            \REG.mem_50_3 , \REG.mem_48_3 , \REG.mem_42_0 , \REG.mem_43_0 , 
            \REG.mem_41_0 , \REG.mem_40_0 , \REG.mem_14_11 , \REG.mem_15_11 , 
            \REG.mem_13_11 , \REG.mem_12_11 , \REG.mem_38_5 , \REG.mem_39_5 , 
            \REG.mem_37_5 , \REG.mem_36_5 , \REG.mem_57_13 , n6121, 
            VCC_net, \fifo_data_out[2] , n6118, \fifo_data_out[1] , 
            \REG.mem_50_1 , \REG.mem_6_9 , \REG.mem_7_9 , \REG.mem_48_1 , 
            n10556, \fifo_data_out[3] , n10562, \fifo_data_out[4] , 
            \REG.mem_18_11 , \REG.mem_16_11 , \REG.mem_5_9 , \REG.mem_4_9 , 
            n10564, \fifo_data_out[5] , n10566, \fifo_data_out[6] , 
            n10568, \fifo_data_out[7] , n10570, \fifo_data_out[8] , 
            n10572, \fifo_data_out[9] , n10574, \fifo_data_out[10] , 
            n10576, \fifo_data_out[11] , \REG.mem_31_5 , n6085, \fifo_data_out[0] , 
            \REG.mem_25_12 , \REG.mem_38_13 , \REG.mem_39_13 , n10578, 
            \fifo_data_out[12] , n10580, \fifo_data_out[13] , \rd_addr_r[6] , 
            \REG.mem_6_15 , \REG.mem_7_15 , n6045, n6043, \REG.mem_5_15 , 
            \REG.mem_4_15 , \REG.mem_35_13 , n6024, n6021, \REG.mem_63_15 , 
            n6020, \REG.mem_63_14 , n6019, \REG.mem_63_13 , n6018, 
            n6017, n6016, \REG.mem_63_10 , n6015, \REG.mem_63_9 , 
            n6014, \REG.mem_63_8 , n6013, \REG.mem_63_7 , n6012, n6011, 
            \REG.mem_63_5 , n6010, \REG.mem_63_4 , n6009, \REG.mem_63_3 , 
            n6008, \REG.mem_63_2 , n6007, \REG.mem_63_1 , n6006, \REG.mem_63_0 , 
            \REG.mem_25_6 , \REG.mem_37_13 , \REG.mem_36_13 , \REG.mem_57_4 , 
            \REG.mem_18_7 , \REG.mem_16_7 , \REG.mem_38_15 , \REG.mem_39_15 , 
            \REG.mem_23_11 , \REG.mem_37_15 , \REG.mem_36_15 , \REG.mem_25_11 , 
            \REG.mem_57_12 , \REG.mem_40_14 , \REG.mem_41_14 , n5953, 
            rp_sync1_r, \REG.mem_42_14 , \REG.mem_43_14 , \REG.mem_46_14 , 
            \REG.mem_47_14 , n5952, n5951, n5950, n5949, n5948, 
            n5947, n5946, n5945, \REG.mem_55_9 , \REG.mem_44_14 , 
            \REG.mem_45_14 , \REG.mem_10_7 , \REG.mem_11_7 , n5928, 
            n5927, n5926, n5924, n5923, n5921, \REG.mem_9_7 , \REG.mem_8_7 , 
            \REG.mem_40_4 , \REG.mem_41_4 , \REG.mem_42_4 , \REG.mem_43_4 , 
            \REG.mem_46_4 , \REG.mem_47_4 , \REG.mem_44_4 , \REG.mem_45_4 , 
            n5901, \REG.mem_57_15 , n5900, \REG.mem_57_14 , n5899, 
            n5898, n5897, \REG.mem_57_11 , n5896, \REG.mem_57_10 , 
            n5895, n5894, \REG.mem_57_8 , n5893, \REG.mem_57_7 , n5892, 
            n5891, \REG.mem_57_5 , n5890, n5889, \REG.mem_57_3 , n5888, 
            \REG.mem_57_2 , n5887, \REG.mem_57_1 , \REG.mem_18_1 , \REG.mem_16_1 , 
            n5885, \REG.mem_35_8 , \REG.mem_38_8 , \REG.mem_39_8 , \REG.mem_36_8 , 
            \REG.mem_37_8 , n5864, wp_sync1_r, n5863, n5862, n5861, 
            n5860, n5859, n5858, \REG.mem_55_15 , n5857, \REG.mem_55_14 , 
            n5856, n5855, n5854, \REG.mem_55_11 , n5853, \rd_sig_diff0_w[0] , 
            n5852, n5851, \REG.mem_55_8 , n5850, n5849, \REG.mem_55_6 , 
            n5848, \REG.mem_55_5 , n5847, \REG.mem_55_4 , n5846, \REG.mem_55_3 , 
            n5845, \REG.mem_55_2 , n5844, \REG.mem_55_1 , n5843, \REG.mem_55_0 , 
            n5842, n5841, n5839, n5838, n5837, \REG.mem_16_15 , 
            \REG.mem_18_15 , \REG.mem_23_15 , n5836, \REG.mem_25_4 , 
            \REG.mem_35_2 , \REG.mem_31_4 , \REG.mem_38_2 , \REG.mem_39_2 , 
            \REG.mem_36_2 , \REG.mem_37_2 , \REG.mem_10_15 , \REG.mem_11_15 , 
            \REG.mem_48_2 , \REG.mem_50_2 , \REG.mem_8_4 , \REG.mem_9_4 , 
            \REG.mem_10_4 , \REG.mem_11_4 , n5771, \REG.mem_50_15 , 
            n5770, \REG.mem_50_14 , n5769, \REG.mem_50_13 , n5768, 
            n5767, \REG.mem_50_11 , n5766, n5765, n5764, \REG.mem_50_8 , 
            n5763, n5762, \REG.mem_50_6 , n5761, \REG.mem_50_5 , n5760, 
            \REG.mem_50_4 , n5759, n5758, n5757, \REG.mem_14_4 , \REG.mem_15_4 , 
            n10873, \REG.mem_12_4 , \REG.mem_13_4 , n10582, \fifo_data_out[14] , 
            n10588, \fifo_data_out[15] , n5753, \REG.mem_50_0 , \REG.mem_3_14 , 
            \REG.mem_6_14 , \REG.mem_7_14 , \REG.mem_4_14 , \REG.mem_5_14 , 
            n5736, \REG.mem_48_15 , n5735, \REG.mem_48_14 , n5734, 
            \REG.mem_48_13 , n5733, n5732, \REG.mem_48_11 , n5731, 
            n5730, n5729, \REG.mem_48_8 , n5728, n5727, \REG.mem_48_6 , 
            n5726, \REG.mem_48_5 , n5725, \REG.mem_48_4 , n5724, n10877, 
            \REG.mem_9_15 , \REG.mem_8_15 , \REG.mem_31_7 , n5723, n5722, 
            n5721, \REG.mem_48_0 , n5720, \REG.mem_47_15 , n5719, 
            n5718, \REG.mem_47_13 , n5717, \REG.mem_47_12 , n5716, 
            \REG.mem_47_11 , n5715, \REG.mem_47_10 , n5714, \REG.mem_47_9 , 
            n5713, n5712, \REG.mem_47_7 , n5711, \REG.mem_47_6 , n5710, 
            \REG.mem_47_5 , n5709, n5708, n5707, \REG.mem_47_2 , n5706, 
            n5705, \REG.mem_47_0 , n5704, \REG.mem_46_15 , n5703, 
            \REG.mem_31_12 , n5702, \REG.mem_46_13 , n5701, \REG.mem_46_12 , 
            n5700, \REG.mem_46_11 , n5699, \REG.mem_46_10 , n5698, 
            \REG.mem_46_9 , n5697, n5696, \REG.mem_46_7 , n5695, \REG.mem_46_6 , 
            n5694, \REG.mem_46_5 , n5693, n5692, n5691, \REG.mem_46_2 , 
            n5690, n5689, \REG.mem_46_0 , n5688, \REG.mem_45_15 , 
            n5687, n5686, \REG.mem_45_13 , n5685, \REG.mem_45_12 , 
            n5684, \REG.mem_45_11 , n5683, \REG.mem_45_10 , n5682, 
            \REG.mem_45_9 , n5681, n5680, \REG.mem_45_7 , n5679, \REG.mem_45_6 , 
            n5678, \REG.mem_45_5 , \REG.mem_38_6 , \REG.mem_39_6 , \REG.mem_37_6 , 
            \REG.mem_36_6 , n5677, \REG.mem_31_11 , n5676, \REG.mem_42_5 , 
            \REG.mem_43_5 , n5675, \REG.mem_45_2 , n5674, n5673, \REG.mem_45_0 , 
            n5671, \REG.mem_44_15 , n5670, n5669, \REG.mem_44_13 , 
            n5668, \REG.mem_44_12 , n5666, \REG.mem_44_11 , n5665, 
            \REG.mem_44_10 , n5664, \REG.mem_44_9 , n5662, n5661, 
            \REG.mem_44_7 , n5660, \REG.mem_44_6 , n5659, \REG.mem_44_5 , 
            n5658, n5657, n5656, \REG.mem_44_2 , n5655, n5654, \REG.mem_44_0 , 
            n5653, \REG.mem_43_15 , n5652, n5651, \REG.mem_43_13 , 
            n5650, \REG.mem_43_12 , n5649, \REG.mem_43_11 , n5648, 
            \REG.mem_43_10 , n5647, \REG.mem_43_9 , n5646, n5645, 
            \REG.mem_43_7 , n5644, \REG.mem_43_6 , \REG.mem_41_5 , \REG.mem_40_5 , 
            \REG.mem_23_1 , \rd_addr_p1_w[0] , \REG.mem_35_11 , n5643, 
            n5642, n5641, n5640, \REG.mem_43_2 , n5639, \REG.mem_43_1 , 
            n5638, n5637, \REG.mem_42_15 , n5636, n5635, \REG.mem_42_13 , 
            n5634, \REG.mem_42_12 , n5633, \REG.mem_42_11 , n5632, 
            \REG.mem_42_10 , n5631, \REG.mem_42_9 , n5630, n5629, 
            \REG.mem_42_7 , n4916, \REG.mem_31_6 , \REG.mem_23_2 , \REG.mem_38_11 , 
            \REG.mem_39_11 , \REG.mem_37_11 , \REG.mem_36_11 , n5628, 
            \REG.mem_42_6 , n5627, n5626, n5625, n5624, \REG.mem_42_2 , 
            n5623, \REG.mem_42_1 , n5622, n5621, \REG.mem_41_15 , 
            n5620, n5619, \REG.mem_41_13 , n5618, \REG.mem_41_12 , 
            n5617, \REG.mem_41_11 , n5616, \REG.mem_41_10 , n5615, 
            \REG.mem_41_9 , n5614, n5613, \REG.mem_41_7 , \REG.mem_3_2 , 
            n5612, \REG.mem_41_6 , n5611, n5610, n5609, n5608, \REG.mem_41_2 , 
            n5607, \REG.mem_41_1 , n5606, n5605, \REG.mem_40_15 , 
            n5604, n5603, \REG.mem_40_13 , n5602, \REG.mem_40_12 , 
            n5601, \REG.mem_40_11 , n5600, \REG.mem_40_10 , n5599, 
            \REG.mem_40_9 , n5598, n5597, \REG.mem_40_7 , \REG.mem_25_9 , 
            n4904, n4903, n4901, n4899, n5596, \REG.mem_40_6 , n5595, 
            n5594, n5593, n5592, \REG.mem_40_2 , n5591, \REG.mem_40_1 , 
            n5590, n5589, n5588, \REG.mem_39_14 , n5587, n5586, 
            \REG.mem_39_12 , n5585, n5584, \REG.mem_39_10 , n5583, 
            \REG.mem_39_9 , n5582, n5581, n4898, \REG.mem_14_1 , \REG.mem_15_1 , 
            DEBUG_5_c, \REG.mem_13_1 , \REG.mem_12_1 , \REG.mem_3_3 , 
            n5580, n5579, n5578, \REG.mem_39_4 , n5577, n5576, n5575, 
            \REG.mem_39_1 , n5573, n5572, n5571, \REG.mem_38_14 , 
            n5570, n5569, \REG.mem_38_12 , n5568, n5567, \REG.mem_38_10 , 
            n5566, \REG.mem_38_9 , n5565, n5564, n5563, n5562, n5561, 
            \REG.mem_38_4 , n5560, n5559, n5558, \REG.mem_38_1 , n5556, 
            n5555, n5554, \REG.mem_37_14 , n5553, n5552, \REG.mem_37_12 , 
            n5551, n5550, \REG.mem_37_10 , n5549, \REG.mem_37_9 , 
            \REG.mem_25_13 , \REG.out_raw[15] , \REG.out_raw[14] , \REG.out_raw[13] , 
            \REG.out_raw[12] , \REG.out_raw[11] , n5548, n5547, n5546, 
            n5545, n5544, \REG.mem_37_4 , n5543, n5542, n5541, \REG.mem_37_1 , 
            n5540, \REG.out_raw[10] , \REG.out_raw[9] , \REG.out_raw[8] , 
            \REG.out_raw[7] , \REG.out_raw[6] , \REG.out_raw[5] , \REG.out_raw[4] , 
            \REG.out_raw[3] , \REG.out_raw[2] , \REG.out_raw[1] , n5526, 
            n5525, \REG.mem_36_14 , n5524, n5523, \REG.mem_36_12 , 
            n5522, n5521, \REG.mem_36_10 , n5520, \REG.mem_36_9 , 
            n5519, n5518, n5517, n5516, \rd_sig_diff0_w[2] , n5515, 
            \REG.mem_36_4 , n5514, n5513, n5512, \REG.mem_36_1 , n5511, 
            n5507, n5506, \REG.mem_35_14 , n5505, n5504, \REG.mem_35_12 , 
            n5503, n5502, \REG.mem_35_10 , n5501, \REG.mem_35_9 , 
            n5500, \rd_sig_diff0_w[1] , n5499, \REG.mem_35_7 , n5498, 
            \REG.mem_35_6 , n5497, \REG.mem_35_5 , n5496, \REG.mem_35_4 , 
            n5495, n5494, n5493, \REG.mem_35_1 , n5492, \REG.mem_6_3 , 
            \REG.mem_7_3 , \REG.mem_5_3 , \REG.mem_4_3 , n5441, n5440, 
            \REG.mem_31_14 , n5439, n5438, n5437, \REG.mem_25_1 , 
            n5436, \REG.mem_31_10 , n58, n5435, \REG.mem_31_9 , n5434, 
            \REG.mem_31_8 , n5433, n5432, n5431, n5430, n5429, n5428, 
            n5427, \REG.mem_31_1 , n5426, n26, DEBUG_1_c_c, write_to_dc32_fifo_latched_N_425, 
            n5345, n5344, \REG.mem_25_14 , n5343, n5342, n5341, 
            n5340, \REG.mem_25_10 , n5339, n5338, \REG.mem_25_8 , 
            n5337, n5336, n5335, n5334, n5333, \REG.mem_25_3 , n5332, 
            n5331, n5330, \REG.mem_25_0 , \REG.mem_14_15 , \REG.mem_15_15 , 
            \REG.mem_6_13 , \REG.mem_7_13 , n5306, n5305, \REG.mem_23_14 , 
            n5304, \REG.mem_23_13 , n5303, n5302, n5301, \REG.mem_23_10 , 
            n5300, \REG.mem_23_9 , n5299, n5298, \REG.mem_23_7 , n5297, 
            \REG.mem_23_6 , n5296, \REG.mem_23_5 , n5295, \REG.mem_23_4 , 
            n5294, \REG.mem_23_3 , n5293, n5292, n5290, \REG.mem_23_0 , 
            \rd_grey_sync_r[5] , \REG.mem_5_13 , \REG.mem_4_13 , \rd_grey_sync_r[4] , 
            \rd_grey_sync_r[3] , \rd_grey_sync_r[2] , \rd_grey_sync_r[1] , 
            \REG.mem_13_15 , \REG.mem_12_15 , n51, n19, \wr_addr_nxt_c[1] , 
            \REG.mem_10_0 , \REG.mem_11_0 , \REG.mem_10_3 , \REG.mem_11_3 , 
            n5224, n5223, \REG.mem_18_14 , n5222, \REG.mem_18_13 , 
            n5221, n5220, \REG.mem_9_3 , \REG.mem_8_3 , \REG.mem_9_0 , 
            \REG.mem_8_0 , \REG.mem_10_13 , \REG.mem_11_13 , n52, \REG.mem_9_13 , 
            \REG.mem_8_13 , n20, n5219, \REG.mem_18_10 , n5218, \REG.mem_18_9 , 
            n5217, n5216, n5215, n5214, \REG.mem_18_5 , n5213, \REG.mem_18_4 , 
            n5212, \REG.mem_18_3 , n5211, n5210, n5209, \REG.mem_18_0 , 
            \REG.mem_14_13 , \REG.mem_15_13 , \REG.mem_13_13 , \REG.mem_12_13 , 
            \REG.mem_6_4 , \REG.mem_7_4 , \REG.mem_5_4 , \REG.mem_4_4 , 
            get_next_word, n5188, n5186, \REG.mem_16_14 , n5185, \REG.mem_16_13 , 
            \REG.mem_6_8 , \REG.mem_7_8 , \REG.mem_3_6 , n5184, \REG.mem_5_8 , 
            \REG.mem_4_8 , \REG.mem_6_2 , \REG.mem_7_2 , \REG.mem_5_2 , 
            \REG.mem_4_2 , rd_fifo_en_w, n5183, n5182, \REG.mem_16_10 , 
            n5181, \REG.mem_16_9 , n5180, n5179, n5178, n5177, \REG.mem_16_5 , 
            n5176, \REG.mem_16_4 , \REG.mem_3_12 , n5175, \REG.mem_16_3 , 
            n5174, n5173, n5172, \REG.mem_16_0 , n5169, n5168, n5167, 
            n47, n5166, n15, n5165, n5164, \REG.mem_15_10 , n5163, 
            \REG.mem_15_9 , n5162, n5161, n5160, \REG.mem_15_6 , n5159, 
            n5158, n5157, \REG.mem_15_3 , n5156, \REG.mem_15_2 , n5155, 
            n5154, \REG.mem_15_0 , n5153, n5152, \REG.mem_6_6 , \REG.mem_7_6 , 
            n5151, n5150, n5149, n5148, \REG.mem_14_10 , n5147, 
            \REG.mem_14_9 , n5146, n5145, n5144, \REG.mem_14_6 , \REG.mem_4_6 , 
            \REG.mem_5_6 , n5143, n5142, n5141, \REG.mem_14_3 , n5140, 
            \REG.mem_14_2 , n5139, n5138, \REG.mem_14_0 , n5137, n5136, 
            n5135, n5134, n5133, n5132, \REG.mem_13_10 , \REG.mem_13_9 , 
            \REG.mem_12_9 , n5131, n5130, n5129, n5128, \REG.mem_13_6 , 
            n5127, n5126, n5125, \REG.mem_13_3 , n5124, \REG.mem_13_2 , 
            n5123, \REG.mem_10_8 , \REG.mem_11_8 , n5122, \REG.mem_13_0 , 
            n5121, n5120, n5119, n5118, \REG.mem_3_9 , \REG.mem_9_8 , 
            \REG.mem_8_8 , n5117, \REG.mem_8_6 , \REG.mem_9_6 , n5116, 
            \REG.mem_12_10 , \REG.mem_10_6 , \REG.mem_11_6 , n53, n21, 
            n5115, n5114, n5113, n5112, \REG.mem_12_6 , n50, n5111, 
            n18, \REG.mem_6_12 , \REG.mem_7_12 , n5110, n5109, \REG.mem_12_3 , 
            n5108, \REG.mem_12_2 , \REG.mem_4_12 , \REG.mem_5_12 , \REG.mem_10_2 , 
            \REG.mem_11_2 , n5107, \REG.mem_9_2 , \REG.mem_8_2 , n54, 
            n22, n5106, \REG.mem_12_0 , \rd_addr_nxt_c_6__N_498[3] , 
            n5105, n5104, n5103, n5102, \REG.mem_11_12 , n5101, 
            n5100, \REG.mem_11_10 , n5099, n5098, n5097, n5096, 
            n5095, \REG.mem_11_5 , n5094, n5093, n5092, n5091, \REG.mem_11_1 , 
            n5090, n5089, n5088, \rd_addr_nxt_c_6__N_498[5] , n5087, 
            n5086, \REG.mem_10_12 , n5085, n5084, \REG.mem_10_10 , 
            n5083, n5082, n5081, n5080, n5079, \REG.mem_10_5 , \REG.mem_10_1 , 
            \REG.mem_9_1 , \REG.mem_8_1 , \rd_addr_nxt_c_6__N_498[2] , 
            n56, n24, n5078, n55, n23, n5077, n40, n8, n5076, 
            n5075, n5074, n5073, n5072, n5071, n5070, \REG.mem_9_12 , 
            n5069, n5068, \REG.mem_9_10 , n5067, n5066, n5065, n57, 
            n5064, n25, n5063, \REG.mem_9_5 , n5062, n5061, n5060, 
            n5059, n5057, n5056, n5055, n5054, n5053, \REG.mem_8_12 , 
            n5052, n5051, \REG.mem_8_10 , n5050, n5049, n5048, n5047, 
            n5046, \REG.mem_8_5 , n5045, n5044, n5043, n5042, n5041, 
            n5040, n5039, n5038, n5037, n5036, n5035, \REG.mem_7_10 , 
            n5034, n5033, n5032, \REG.mem_7_7 , n5031, n5030, \REG.mem_7_5 , 
            n5029, n5028, n5027, n5026, n5025, \REG.mem_7_0 , n5024, 
            n5023, n5022, n5021, n5020, n5019, \REG.mem_6_10 , n5018, 
            n5017, n5016, \REG.mem_6_7 , n5015, n5014, \REG.mem_6_5 , 
            n5013, n5012, n5011, n5010, n5009, \REG.mem_6_0 , n5008, 
            n5007, n5006, n5005, n5004, n5003, \REG.mem_5_10 , n5002, 
            n5001, n5000, \REG.mem_5_7 , n4999, n4998, \REG.mem_5_5 , 
            n4997, n4996, n4995, n4994, n4993, \REG.mem_5_0 , n4992, 
            n4991, n4990, n4989, n4988, n4987, \REG.mem_4_10 , n4986, 
            n4985, n4984, \REG.mem_4_7 , n4983, n4982, \REG.mem_4_5 , 
            n4981, n4980, n4979, n4978, n4977, \REG.mem_4_0 , n4976, 
            n4975, n4974, n4973, n4972, n4971, \REG.mem_3_10 , n4970, 
            n4969, \REG.mem_3_8 , FT_OE_N_420, n49, n17, n42, n10, 
            n4968, \REG.mem_3_7 , n4967, n4966, \REG.mem_3_5 , n4965, 
            n34, n4964, n4963, n2, n4962, n4961, \REG.mem_3_0 , 
            n59, n27, n60, n28, n61, n29) /* synthesis syn_module_defined=1 */ ;
    output \rd_addr_r[0] ;
    output \REG.mem_14_5 ;
    output \REG.mem_15_5 ;
    input \dc32_fifo_data_in[6] ;
    output dc32_fifo_almost_full;
    input FIFO_CLK_c;
    input reset_per_frame;
    output \REG.mem_13_5 ;
    output \REG.mem_12_5 ;
    input \dc32_fifo_data_in[5] ;
    input \dc32_fifo_data_in[4] ;
    output \REG.mem_31_0 ;
    input GND_net;
    input \dc32_fifo_data_in[3] ;
    output \REG.mem_55_13 ;
    input \dc32_fifo_data_in[2] ;
    output \REG.mem_38_7 ;
    output \REG.mem_39_7 ;
    output \REG.mem_36_7 ;
    output \REG.mem_37_7 ;
    output \REG.mem_16_8 ;
    output \REG.mem_18_8 ;
    output \REG.mem_3_13 ;
    output \REG.mem_57_6 ;
    input \dc32_fifo_data_in[1] ;
    output \REG.mem_63_11 ;
    input \dc32_fifo_data_in[0] ;
    output \REG.mem_35_0 ;
    output t_rd_fifo_en_w;
    output \REG.out_raw[0] ;
    input SLM_CLK_c;
    output \REG.mem_55_10 ;
    output n62;
    output n30;
    output \REG.mem_31_3 ;
    output \REG.mem_48_7 ;
    output \REG.mem_50_7 ;
    output \REG.mem_55_7 ;
    output \REG.mem_48_10 ;
    output \REG.mem_50_10 ;
    output [6:0]wr_grey_sync_r;
    output \wr_addr_nxt_c[5] ;
    output \REG.mem_23_8 ;
    output \REG.mem_25_5 ;
    output \rd_grey_sync_r[0] ;
    output \REG.mem_25_15 ;
    output \REG.mem_14_12 ;
    output \REG.mem_15_12 ;
    output DEBUG_3_c;
    output \REG.mem_13_12 ;
    output \REG.mem_12_12 ;
    input \aempty_flag_impl.ae_flag_nxt_w ;
    output dc32_fifo_almost_empty;
    output \REG.mem_6_1 ;
    output \REG.mem_7_1 ;
    output \REG.mem_5_1 ;
    output \REG.mem_4_1 ;
    output \REG.mem_57_9 ;
    output \REG.mem_35_3 ;
    output \REG.mem_46_1 ;
    output \REG.mem_47_1 ;
    output \REG.mem_45_1 ;
    output \REG.mem_44_1 ;
    output \REG.mem_25_2 ;
    input \dc32_fifo_data_in[15] ;
    input \dc32_fifo_data_in[14] ;
    input \dc32_fifo_data_in[13] ;
    output \REG.mem_3_11 ;
    output \REG.mem_31_2 ;
    output \REG.mem_50_12 ;
    input \dc32_fifo_data_in[12] ;
    output \REG.mem_6_11 ;
    output \REG.mem_7_11 ;
    output \REG.mem_5_11 ;
    output \REG.mem_4_11 ;
    input \dc32_fifo_data_in[11] ;
    output \REG.mem_48_12 ;
    output \REG.mem_3_4 ;
    output \REG.mem_14_8 ;
    output \REG.mem_15_8 ;
    output \REG.mem_8_14 ;
    output \REG.mem_9_14 ;
    input \dc32_fifo_data_in[10] ;
    output \REG.mem_10_14 ;
    output \REG.mem_11_14 ;
    output \REG.mem_63_6 ;
    output \REG.mem_13_8 ;
    output \REG.mem_12_8 ;
    output \REG.mem_14_14 ;
    output \REG.mem_15_14 ;
    input \dc32_fifo_data_in[9] ;
    input \dc32_fifo_data_in[8] ;
    output \REG.mem_3_1 ;
    input \dc32_fifo_data_in[7] ;
    output \REG.mem_12_14 ;
    output \REG.mem_13_14 ;
    output \REG.mem_42_8 ;
    output \REG.mem_43_8 ;
    output \REG.mem_41_8 ;
    output \REG.mem_40_8 ;
    output \REG.mem_18_12 ;
    output \REG.mem_16_12 ;
    output \REG.mem_31_15 ;
    output \REG.mem_38_3 ;
    output \REG.mem_39_3 ;
    output \REG.mem_37_3 ;
    output \REG.mem_36_3 ;
    output \REG.mem_42_3 ;
    output \REG.mem_43_3 ;
    output \REG.mem_14_7 ;
    output \REG.mem_15_7 ;
    output \REG.mem_13_7 ;
    output \REG.mem_12_7 ;
    output \REG.mem_41_3 ;
    output \REG.mem_40_3 ;
    output \REG.mem_57_0 ;
    output \REG.mem_10_11 ;
    output \REG.mem_11_11 ;
    output \REG.mem_9_11 ;
    output \REG.mem_8_11 ;
    output \REG.mem_63_12 ;
    output \REG.mem_55_12 ;
    output \REG.mem_35_15 ;
    output \REG.mem_3_15 ;
    output \wr_addr_nxt_c[3] ;
    output \REG.mem_50_9 ;
    output \REG.mem_48_9 ;
    output \REG.mem_46_8 ;
    output \REG.mem_47_8 ;
    output \REG.mem_46_3 ;
    output \REG.mem_47_3 ;
    output \REG.mem_45_8 ;
    output \REG.mem_44_8 ;
    output \REG.mem_16_2 ;
    output \REG.mem_10_9 ;
    output \REG.mem_11_9 ;
    output \REG.mem_45_3 ;
    output \REG.mem_44_3 ;
    output \REG.mem_25_7 ;
    output \REG.mem_23_12 ;
    output \REG.mem_18_2 ;
    output \REG.mem_38_0 ;
    output \REG.mem_39_0 ;
    output \REG.mem_31_13 ;
    output \REG.mem_37_0 ;
    output \REG.mem_36_0 ;
    output \REG.mem_18_6 ;
    output \REG.mem_16_6 ;
    output \REG.mem_9_9 ;
    output \REG.mem_8_9 ;
    output \REG.mem_50_3 ;
    output \REG.mem_48_3 ;
    output \REG.mem_42_0 ;
    output \REG.mem_43_0 ;
    output \REG.mem_41_0 ;
    output \REG.mem_40_0 ;
    output \REG.mem_14_11 ;
    output \REG.mem_15_11 ;
    output \REG.mem_13_11 ;
    output \REG.mem_12_11 ;
    output \REG.mem_38_5 ;
    output \REG.mem_39_5 ;
    output \REG.mem_37_5 ;
    output \REG.mem_36_5 ;
    output \REG.mem_57_13 ;
    input n6121;
    input VCC_net;
    output \fifo_data_out[2] ;
    input n6118;
    output \fifo_data_out[1] ;
    output \REG.mem_50_1 ;
    output \REG.mem_6_9 ;
    output \REG.mem_7_9 ;
    output \REG.mem_48_1 ;
    input n10556;
    output \fifo_data_out[3] ;
    input n10562;
    output \fifo_data_out[4] ;
    output \REG.mem_18_11 ;
    output \REG.mem_16_11 ;
    output \REG.mem_5_9 ;
    output \REG.mem_4_9 ;
    input n10564;
    output \fifo_data_out[5] ;
    input n10566;
    output \fifo_data_out[6] ;
    input n10568;
    output \fifo_data_out[7] ;
    input n10570;
    output \fifo_data_out[8] ;
    input n10572;
    output \fifo_data_out[9] ;
    input n10574;
    output \fifo_data_out[10] ;
    input n10576;
    output \fifo_data_out[11] ;
    output \REG.mem_31_5 ;
    input n6085;
    output \fifo_data_out[0] ;
    output \REG.mem_25_12 ;
    output \REG.mem_38_13 ;
    output \REG.mem_39_13 ;
    input n10578;
    output \fifo_data_out[12] ;
    input n10580;
    output \fifo_data_out[13] ;
    output \rd_addr_r[6] ;
    output \REG.mem_6_15 ;
    output \REG.mem_7_15 ;
    input n6045;
    input n6043;
    output \REG.mem_5_15 ;
    output \REG.mem_4_15 ;
    output \REG.mem_35_13 ;
    input n6024;
    input n6021;
    output \REG.mem_63_15 ;
    input n6020;
    output \REG.mem_63_14 ;
    input n6019;
    output \REG.mem_63_13 ;
    input n6018;
    input n6017;
    input n6016;
    output \REG.mem_63_10 ;
    input n6015;
    output \REG.mem_63_9 ;
    input n6014;
    output \REG.mem_63_8 ;
    input n6013;
    output \REG.mem_63_7 ;
    input n6012;
    input n6011;
    output \REG.mem_63_5 ;
    input n6010;
    output \REG.mem_63_4 ;
    input n6009;
    output \REG.mem_63_3 ;
    input n6008;
    output \REG.mem_63_2 ;
    input n6007;
    output \REG.mem_63_1 ;
    input n6006;
    output \REG.mem_63_0 ;
    output \REG.mem_25_6 ;
    output \REG.mem_37_13 ;
    output \REG.mem_36_13 ;
    output \REG.mem_57_4 ;
    output \REG.mem_18_7 ;
    output \REG.mem_16_7 ;
    output \REG.mem_38_15 ;
    output \REG.mem_39_15 ;
    output \REG.mem_23_11 ;
    output \REG.mem_37_15 ;
    output \REG.mem_36_15 ;
    output \REG.mem_25_11 ;
    output \REG.mem_57_12 ;
    output \REG.mem_40_14 ;
    output \REG.mem_41_14 ;
    input n5953;
    output [6:0]rp_sync1_r;
    output \REG.mem_42_14 ;
    output \REG.mem_43_14 ;
    output \REG.mem_46_14 ;
    output \REG.mem_47_14 ;
    input n5952;
    input n5951;
    input n5950;
    input n5949;
    input n5948;
    input n5947;
    input n5946;
    input n5945;
    output \REG.mem_55_9 ;
    output \REG.mem_44_14 ;
    output \REG.mem_45_14 ;
    output \REG.mem_10_7 ;
    output \REG.mem_11_7 ;
    input n5928;
    input n5927;
    input n5926;
    input n5924;
    input n5923;
    input n5921;
    output \REG.mem_9_7 ;
    output \REG.mem_8_7 ;
    output \REG.mem_40_4 ;
    output \REG.mem_41_4 ;
    output \REG.mem_42_4 ;
    output \REG.mem_43_4 ;
    output \REG.mem_46_4 ;
    output \REG.mem_47_4 ;
    output \REG.mem_44_4 ;
    output \REG.mem_45_4 ;
    input n5901;
    output \REG.mem_57_15 ;
    input n5900;
    output \REG.mem_57_14 ;
    input n5899;
    input n5898;
    input n5897;
    output \REG.mem_57_11 ;
    input n5896;
    output \REG.mem_57_10 ;
    input n5895;
    input n5894;
    output \REG.mem_57_8 ;
    input n5893;
    output \REG.mem_57_7 ;
    input n5892;
    input n5891;
    output \REG.mem_57_5 ;
    input n5890;
    input n5889;
    output \REG.mem_57_3 ;
    input n5888;
    output \REG.mem_57_2 ;
    input n5887;
    output \REG.mem_57_1 ;
    output \REG.mem_18_1 ;
    output \REG.mem_16_1 ;
    input n5885;
    output \REG.mem_35_8 ;
    output \REG.mem_38_8 ;
    output \REG.mem_39_8 ;
    output \REG.mem_36_8 ;
    output \REG.mem_37_8 ;
    input n5864;
    output [6:0]wp_sync1_r;
    input n5863;
    input n5862;
    input n5861;
    input n5860;
    input n5859;
    input n5858;
    output \REG.mem_55_15 ;
    input n5857;
    output \REG.mem_55_14 ;
    input n5856;
    input n5855;
    input n5854;
    output \REG.mem_55_11 ;
    input n5853;
    output \rd_sig_diff0_w[0] ;
    input n5852;
    input n5851;
    output \REG.mem_55_8 ;
    input n5850;
    input n5849;
    output \REG.mem_55_6 ;
    input n5848;
    output \REG.mem_55_5 ;
    input n5847;
    output \REG.mem_55_4 ;
    input n5846;
    output \REG.mem_55_3 ;
    input n5845;
    output \REG.mem_55_2 ;
    input n5844;
    output \REG.mem_55_1 ;
    input n5843;
    output \REG.mem_55_0 ;
    input n5842;
    input n5841;
    input n5839;
    input n5838;
    input n5837;
    output \REG.mem_16_15 ;
    output \REG.mem_18_15 ;
    output \REG.mem_23_15 ;
    input n5836;
    output \REG.mem_25_4 ;
    output \REG.mem_35_2 ;
    output \REG.mem_31_4 ;
    output \REG.mem_38_2 ;
    output \REG.mem_39_2 ;
    output \REG.mem_36_2 ;
    output \REG.mem_37_2 ;
    output \REG.mem_10_15 ;
    output \REG.mem_11_15 ;
    output \REG.mem_48_2 ;
    output \REG.mem_50_2 ;
    output \REG.mem_8_4 ;
    output \REG.mem_9_4 ;
    output \REG.mem_10_4 ;
    output \REG.mem_11_4 ;
    input n5771;
    output \REG.mem_50_15 ;
    input n5770;
    output \REG.mem_50_14 ;
    input n5769;
    output \REG.mem_50_13 ;
    input n5768;
    input n5767;
    output \REG.mem_50_11 ;
    input n5766;
    input n5765;
    input n5764;
    output \REG.mem_50_8 ;
    input n5763;
    input n5762;
    output \REG.mem_50_6 ;
    input n5761;
    output \REG.mem_50_5 ;
    input n5760;
    output \REG.mem_50_4 ;
    input n5759;
    input n5758;
    input n5757;
    output \REG.mem_14_4 ;
    output \REG.mem_15_4 ;
    output n10873;
    output \REG.mem_12_4 ;
    output \REG.mem_13_4 ;
    input n10582;
    output \fifo_data_out[14] ;
    input n10588;
    output \fifo_data_out[15] ;
    input n5753;
    output \REG.mem_50_0 ;
    output \REG.mem_3_14 ;
    output \REG.mem_6_14 ;
    output \REG.mem_7_14 ;
    output \REG.mem_4_14 ;
    output \REG.mem_5_14 ;
    input n5736;
    output \REG.mem_48_15 ;
    input n5735;
    output \REG.mem_48_14 ;
    input n5734;
    output \REG.mem_48_13 ;
    input n5733;
    input n5732;
    output \REG.mem_48_11 ;
    input n5731;
    input n5730;
    input n5729;
    output \REG.mem_48_8 ;
    input n5728;
    input n5727;
    output \REG.mem_48_6 ;
    input n5726;
    output \REG.mem_48_5 ;
    input n5725;
    output \REG.mem_48_4 ;
    input n5724;
    output n10877;
    output \REG.mem_9_15 ;
    output \REG.mem_8_15 ;
    output \REG.mem_31_7 ;
    input n5723;
    input n5722;
    input n5721;
    output \REG.mem_48_0 ;
    input n5720;
    output \REG.mem_47_15 ;
    input n5719;
    input n5718;
    output \REG.mem_47_13 ;
    input n5717;
    output \REG.mem_47_12 ;
    input n5716;
    output \REG.mem_47_11 ;
    input n5715;
    output \REG.mem_47_10 ;
    input n5714;
    output \REG.mem_47_9 ;
    input n5713;
    input n5712;
    output \REG.mem_47_7 ;
    input n5711;
    output \REG.mem_47_6 ;
    input n5710;
    output \REG.mem_47_5 ;
    input n5709;
    input n5708;
    input n5707;
    output \REG.mem_47_2 ;
    input n5706;
    input n5705;
    output \REG.mem_47_0 ;
    input n5704;
    output \REG.mem_46_15 ;
    input n5703;
    output \REG.mem_31_12 ;
    input n5702;
    output \REG.mem_46_13 ;
    input n5701;
    output \REG.mem_46_12 ;
    input n5700;
    output \REG.mem_46_11 ;
    input n5699;
    output \REG.mem_46_10 ;
    input n5698;
    output \REG.mem_46_9 ;
    input n5697;
    input n5696;
    output \REG.mem_46_7 ;
    input n5695;
    output \REG.mem_46_6 ;
    input n5694;
    output \REG.mem_46_5 ;
    input n5693;
    input n5692;
    input n5691;
    output \REG.mem_46_2 ;
    input n5690;
    input n5689;
    output \REG.mem_46_0 ;
    input n5688;
    output \REG.mem_45_15 ;
    input n5687;
    input n5686;
    output \REG.mem_45_13 ;
    input n5685;
    output \REG.mem_45_12 ;
    input n5684;
    output \REG.mem_45_11 ;
    input n5683;
    output \REG.mem_45_10 ;
    input n5682;
    output \REG.mem_45_9 ;
    input n5681;
    input n5680;
    output \REG.mem_45_7 ;
    input n5679;
    output \REG.mem_45_6 ;
    input n5678;
    output \REG.mem_45_5 ;
    output \REG.mem_38_6 ;
    output \REG.mem_39_6 ;
    output \REG.mem_37_6 ;
    output \REG.mem_36_6 ;
    input n5677;
    output \REG.mem_31_11 ;
    input n5676;
    output \REG.mem_42_5 ;
    output \REG.mem_43_5 ;
    input n5675;
    output \REG.mem_45_2 ;
    input n5674;
    input n5673;
    output \REG.mem_45_0 ;
    input n5671;
    output \REG.mem_44_15 ;
    input n5670;
    input n5669;
    output \REG.mem_44_13 ;
    input n5668;
    output \REG.mem_44_12 ;
    input n5666;
    output \REG.mem_44_11 ;
    input n5665;
    output \REG.mem_44_10 ;
    input n5664;
    output \REG.mem_44_9 ;
    input n5662;
    input n5661;
    output \REG.mem_44_7 ;
    input n5660;
    output \REG.mem_44_6 ;
    input n5659;
    output \REG.mem_44_5 ;
    input n5658;
    input n5657;
    input n5656;
    output \REG.mem_44_2 ;
    input n5655;
    input n5654;
    output \REG.mem_44_0 ;
    input n5653;
    output \REG.mem_43_15 ;
    input n5652;
    input n5651;
    output \REG.mem_43_13 ;
    input n5650;
    output \REG.mem_43_12 ;
    input n5649;
    output \REG.mem_43_11 ;
    input n5648;
    output \REG.mem_43_10 ;
    input n5647;
    output \REG.mem_43_9 ;
    input n5646;
    input n5645;
    output \REG.mem_43_7 ;
    input n5644;
    output \REG.mem_43_6 ;
    output \REG.mem_41_5 ;
    output \REG.mem_40_5 ;
    output \REG.mem_23_1 ;
    output \rd_addr_p1_w[0] ;
    output \REG.mem_35_11 ;
    input n5643;
    input n5642;
    input n5641;
    input n5640;
    output \REG.mem_43_2 ;
    input n5639;
    output \REG.mem_43_1 ;
    input n5638;
    input n5637;
    output \REG.mem_42_15 ;
    input n5636;
    input n5635;
    output \REG.mem_42_13 ;
    input n5634;
    output \REG.mem_42_12 ;
    input n5633;
    output \REG.mem_42_11 ;
    input n5632;
    output \REG.mem_42_10 ;
    input n5631;
    output \REG.mem_42_9 ;
    input n5630;
    input n5629;
    output \REG.mem_42_7 ;
    input n4916;
    output \REG.mem_31_6 ;
    output \REG.mem_23_2 ;
    output \REG.mem_38_11 ;
    output \REG.mem_39_11 ;
    output \REG.mem_37_11 ;
    output \REG.mem_36_11 ;
    input n5628;
    output \REG.mem_42_6 ;
    input n5627;
    input n5626;
    input n5625;
    input n5624;
    output \REG.mem_42_2 ;
    input n5623;
    output \REG.mem_42_1 ;
    input n5622;
    input n5621;
    output \REG.mem_41_15 ;
    input n5620;
    input n5619;
    output \REG.mem_41_13 ;
    input n5618;
    output \REG.mem_41_12 ;
    input n5617;
    output \REG.mem_41_11 ;
    input n5616;
    output \REG.mem_41_10 ;
    input n5615;
    output \REG.mem_41_9 ;
    input n5614;
    input n5613;
    output \REG.mem_41_7 ;
    output \REG.mem_3_2 ;
    input n5612;
    output \REG.mem_41_6 ;
    input n5611;
    input n5610;
    input n5609;
    input n5608;
    output \REG.mem_41_2 ;
    input n5607;
    output \REG.mem_41_1 ;
    input n5606;
    input n5605;
    output \REG.mem_40_15 ;
    input n5604;
    input n5603;
    output \REG.mem_40_13 ;
    input n5602;
    output \REG.mem_40_12 ;
    input n5601;
    output \REG.mem_40_11 ;
    input n5600;
    output \REG.mem_40_10 ;
    input n5599;
    output \REG.mem_40_9 ;
    input n5598;
    input n5597;
    output \REG.mem_40_7 ;
    output \REG.mem_25_9 ;
    input n4904;
    input n4903;
    input n4901;
    input n4899;
    input n5596;
    output \REG.mem_40_6 ;
    input n5595;
    input n5594;
    input n5593;
    input n5592;
    output \REG.mem_40_2 ;
    input n5591;
    output \REG.mem_40_1 ;
    input n5590;
    input n5589;
    input n5588;
    output \REG.mem_39_14 ;
    input n5587;
    input n5586;
    output \REG.mem_39_12 ;
    input n5585;
    input n5584;
    output \REG.mem_39_10 ;
    input n5583;
    output \REG.mem_39_9 ;
    input n5582;
    input n5581;
    input n4898;
    output \REG.mem_14_1 ;
    output \REG.mem_15_1 ;
    input DEBUG_5_c;
    output \REG.mem_13_1 ;
    output \REG.mem_12_1 ;
    output \REG.mem_3_3 ;
    input n5580;
    input n5579;
    input n5578;
    output \REG.mem_39_4 ;
    input n5577;
    input n5576;
    input n5575;
    output \REG.mem_39_1 ;
    input n5573;
    input n5572;
    input n5571;
    output \REG.mem_38_14 ;
    input n5570;
    input n5569;
    output \REG.mem_38_12 ;
    input n5568;
    input n5567;
    output \REG.mem_38_10 ;
    input n5566;
    output \REG.mem_38_9 ;
    input n5565;
    input n5564;
    input n5563;
    input n5562;
    input n5561;
    output \REG.mem_38_4 ;
    input n5560;
    input n5559;
    input n5558;
    output \REG.mem_38_1 ;
    input n5556;
    input n5555;
    input n5554;
    output \REG.mem_37_14 ;
    input n5553;
    input n5552;
    output \REG.mem_37_12 ;
    input n5551;
    input n5550;
    output \REG.mem_37_10 ;
    input n5549;
    output \REG.mem_37_9 ;
    output \REG.mem_25_13 ;
    output \REG.out_raw[15] ;
    output \REG.out_raw[14] ;
    output \REG.out_raw[13] ;
    output \REG.out_raw[12] ;
    output \REG.out_raw[11] ;
    input n5548;
    input n5547;
    input n5546;
    input n5545;
    input n5544;
    output \REG.mem_37_4 ;
    input n5543;
    input n5542;
    input n5541;
    output \REG.mem_37_1 ;
    input n5540;
    output \REG.out_raw[10] ;
    output \REG.out_raw[9] ;
    output \REG.out_raw[8] ;
    output \REG.out_raw[7] ;
    output \REG.out_raw[6] ;
    output \REG.out_raw[5] ;
    output \REG.out_raw[4] ;
    output \REG.out_raw[3] ;
    output \REG.out_raw[2] ;
    output \REG.out_raw[1] ;
    input n5526;
    input n5525;
    output \REG.mem_36_14 ;
    input n5524;
    input n5523;
    output \REG.mem_36_12 ;
    input n5522;
    input n5521;
    output \REG.mem_36_10 ;
    input n5520;
    output \REG.mem_36_9 ;
    input n5519;
    input n5518;
    input n5517;
    input n5516;
    output \rd_sig_diff0_w[2] ;
    input n5515;
    output \REG.mem_36_4 ;
    input n5514;
    input n5513;
    input n5512;
    output \REG.mem_36_1 ;
    input n5511;
    input n5507;
    input n5506;
    output \REG.mem_35_14 ;
    input n5505;
    input n5504;
    output \REG.mem_35_12 ;
    input n5503;
    input n5502;
    output \REG.mem_35_10 ;
    input n5501;
    output \REG.mem_35_9 ;
    input n5500;
    output \rd_sig_diff0_w[1] ;
    input n5499;
    output \REG.mem_35_7 ;
    input n5498;
    output \REG.mem_35_6 ;
    input n5497;
    output \REG.mem_35_5 ;
    input n5496;
    output \REG.mem_35_4 ;
    input n5495;
    input n5494;
    input n5493;
    output \REG.mem_35_1 ;
    input n5492;
    output \REG.mem_6_3 ;
    output \REG.mem_7_3 ;
    output \REG.mem_5_3 ;
    output \REG.mem_4_3 ;
    input n5441;
    input n5440;
    output \REG.mem_31_14 ;
    input n5439;
    input n5438;
    input n5437;
    output \REG.mem_25_1 ;
    input n5436;
    output \REG.mem_31_10 ;
    output n58;
    input n5435;
    output \REG.mem_31_9 ;
    input n5434;
    output \REG.mem_31_8 ;
    input n5433;
    input n5432;
    input n5431;
    input n5430;
    input n5429;
    input n5428;
    input n5427;
    output \REG.mem_31_1 ;
    input n5426;
    output n26;
    input DEBUG_1_c_c;
    output write_to_dc32_fifo_latched_N_425;
    input n5345;
    input n5344;
    output \REG.mem_25_14 ;
    input n5343;
    input n5342;
    input n5341;
    input n5340;
    output \REG.mem_25_10 ;
    input n5339;
    input n5338;
    output \REG.mem_25_8 ;
    input n5337;
    input n5336;
    input n5335;
    input n5334;
    input n5333;
    output \REG.mem_25_3 ;
    input n5332;
    input n5331;
    input n5330;
    output \REG.mem_25_0 ;
    output \REG.mem_14_15 ;
    output \REG.mem_15_15 ;
    output \REG.mem_6_13 ;
    output \REG.mem_7_13 ;
    input n5306;
    input n5305;
    output \REG.mem_23_14 ;
    input n5304;
    output \REG.mem_23_13 ;
    input n5303;
    input n5302;
    input n5301;
    output \REG.mem_23_10 ;
    input n5300;
    output \REG.mem_23_9 ;
    input n5299;
    input n5298;
    output \REG.mem_23_7 ;
    input n5297;
    output \REG.mem_23_6 ;
    input n5296;
    output \REG.mem_23_5 ;
    input n5295;
    output \REG.mem_23_4 ;
    input n5294;
    output \REG.mem_23_3 ;
    input n5293;
    input n5292;
    input n5290;
    output \REG.mem_23_0 ;
    output \rd_grey_sync_r[5] ;
    output \REG.mem_5_13 ;
    output \REG.mem_4_13 ;
    output \rd_grey_sync_r[4] ;
    output \rd_grey_sync_r[3] ;
    output \rd_grey_sync_r[2] ;
    output \rd_grey_sync_r[1] ;
    output \REG.mem_13_15 ;
    output \REG.mem_12_15 ;
    output n51;
    output n19;
    output \wr_addr_nxt_c[1] ;
    output \REG.mem_10_0 ;
    output \REG.mem_11_0 ;
    output \REG.mem_10_3 ;
    output \REG.mem_11_3 ;
    input n5224;
    input n5223;
    output \REG.mem_18_14 ;
    input n5222;
    output \REG.mem_18_13 ;
    input n5221;
    input n5220;
    output \REG.mem_9_3 ;
    output \REG.mem_8_3 ;
    output \REG.mem_9_0 ;
    output \REG.mem_8_0 ;
    output \REG.mem_10_13 ;
    output \REG.mem_11_13 ;
    output n52;
    output \REG.mem_9_13 ;
    output \REG.mem_8_13 ;
    output n20;
    input n5219;
    output \REG.mem_18_10 ;
    input n5218;
    output \REG.mem_18_9 ;
    input n5217;
    input n5216;
    input n5215;
    input n5214;
    output \REG.mem_18_5 ;
    input n5213;
    output \REG.mem_18_4 ;
    input n5212;
    output \REG.mem_18_3 ;
    input n5211;
    input n5210;
    input n5209;
    output \REG.mem_18_0 ;
    output \REG.mem_14_13 ;
    output \REG.mem_15_13 ;
    output \REG.mem_13_13 ;
    output \REG.mem_12_13 ;
    output \REG.mem_6_4 ;
    output \REG.mem_7_4 ;
    output \REG.mem_5_4 ;
    output \REG.mem_4_4 ;
    input get_next_word;
    input n5188;
    input n5186;
    output \REG.mem_16_14 ;
    input n5185;
    output \REG.mem_16_13 ;
    output \REG.mem_6_8 ;
    output \REG.mem_7_8 ;
    output \REG.mem_3_6 ;
    input n5184;
    output \REG.mem_5_8 ;
    output \REG.mem_4_8 ;
    output \REG.mem_6_2 ;
    output \REG.mem_7_2 ;
    output \REG.mem_5_2 ;
    output \REG.mem_4_2 ;
    output rd_fifo_en_w;
    input n5183;
    input n5182;
    output \REG.mem_16_10 ;
    input n5181;
    output \REG.mem_16_9 ;
    input n5180;
    input n5179;
    input n5178;
    input n5177;
    output \REG.mem_16_5 ;
    input n5176;
    output \REG.mem_16_4 ;
    output \REG.mem_3_12 ;
    input n5175;
    output \REG.mem_16_3 ;
    input n5174;
    input n5173;
    input n5172;
    output \REG.mem_16_0 ;
    input n5169;
    input n5168;
    input n5167;
    output n47;
    input n5166;
    output n15;
    input n5165;
    input n5164;
    output \REG.mem_15_10 ;
    input n5163;
    output \REG.mem_15_9 ;
    input n5162;
    input n5161;
    input n5160;
    output \REG.mem_15_6 ;
    input n5159;
    input n5158;
    input n5157;
    output \REG.mem_15_3 ;
    input n5156;
    output \REG.mem_15_2 ;
    input n5155;
    input n5154;
    output \REG.mem_15_0 ;
    input n5153;
    input n5152;
    output \REG.mem_6_6 ;
    output \REG.mem_7_6 ;
    input n5151;
    input n5150;
    input n5149;
    input n5148;
    output \REG.mem_14_10 ;
    input n5147;
    output \REG.mem_14_9 ;
    input n5146;
    input n5145;
    input n5144;
    output \REG.mem_14_6 ;
    output \REG.mem_4_6 ;
    output \REG.mem_5_6 ;
    input n5143;
    input n5142;
    input n5141;
    output \REG.mem_14_3 ;
    input n5140;
    output \REG.mem_14_2 ;
    input n5139;
    input n5138;
    output \REG.mem_14_0 ;
    input n5137;
    input n5136;
    input n5135;
    input n5134;
    input n5133;
    input n5132;
    output \REG.mem_13_10 ;
    output \REG.mem_13_9 ;
    output \REG.mem_12_9 ;
    input n5131;
    input n5130;
    input n5129;
    input n5128;
    output \REG.mem_13_6 ;
    input n5127;
    input n5126;
    input n5125;
    output \REG.mem_13_3 ;
    input n5124;
    output \REG.mem_13_2 ;
    input n5123;
    output \REG.mem_10_8 ;
    output \REG.mem_11_8 ;
    input n5122;
    output \REG.mem_13_0 ;
    input n5121;
    input n5120;
    input n5119;
    input n5118;
    output \REG.mem_3_9 ;
    output \REG.mem_9_8 ;
    output \REG.mem_8_8 ;
    input n5117;
    output \REG.mem_8_6 ;
    output \REG.mem_9_6 ;
    input n5116;
    output \REG.mem_12_10 ;
    output \REG.mem_10_6 ;
    output \REG.mem_11_6 ;
    output n53;
    output n21;
    input n5115;
    input n5114;
    input n5113;
    input n5112;
    output \REG.mem_12_6 ;
    output n50;
    input n5111;
    output n18;
    output \REG.mem_6_12 ;
    output \REG.mem_7_12 ;
    input n5110;
    input n5109;
    output \REG.mem_12_3 ;
    input n5108;
    output \REG.mem_12_2 ;
    output \REG.mem_4_12 ;
    output \REG.mem_5_12 ;
    output \REG.mem_10_2 ;
    output \REG.mem_11_2 ;
    input n5107;
    output \REG.mem_9_2 ;
    output \REG.mem_8_2 ;
    output n54;
    output n22;
    input n5106;
    output \REG.mem_12_0 ;
    output \rd_addr_nxt_c_6__N_498[3] ;
    input n5105;
    input n5104;
    input n5103;
    input n5102;
    output \REG.mem_11_12 ;
    input n5101;
    input n5100;
    output \REG.mem_11_10 ;
    input n5099;
    input n5098;
    input n5097;
    input n5096;
    input n5095;
    output \REG.mem_11_5 ;
    input n5094;
    input n5093;
    input n5092;
    input n5091;
    output \REG.mem_11_1 ;
    input n5090;
    input n5089;
    input n5088;
    output \rd_addr_nxt_c_6__N_498[5] ;
    input n5087;
    input n5086;
    output \REG.mem_10_12 ;
    input n5085;
    input n5084;
    output \REG.mem_10_10 ;
    input n5083;
    input n5082;
    input n5081;
    input n5080;
    input n5079;
    output \REG.mem_10_5 ;
    output \REG.mem_10_1 ;
    output \REG.mem_9_1 ;
    output \REG.mem_8_1 ;
    output \rd_addr_nxt_c_6__N_498[2] ;
    output n56;
    output n24;
    input n5078;
    output n55;
    output n23;
    input n5077;
    output n40;
    output n8;
    input n5076;
    input n5075;
    input n5074;
    input n5073;
    input n5072;
    input n5071;
    input n5070;
    output \REG.mem_9_12 ;
    input n5069;
    input n5068;
    output \REG.mem_9_10 ;
    input n5067;
    input n5066;
    input n5065;
    output n57;
    input n5064;
    output n25;
    input n5063;
    output \REG.mem_9_5 ;
    input n5062;
    input n5061;
    input n5060;
    input n5059;
    input n5057;
    input n5056;
    input n5055;
    input n5054;
    input n5053;
    output \REG.mem_8_12 ;
    input n5052;
    input n5051;
    output \REG.mem_8_10 ;
    input n5050;
    input n5049;
    input n5048;
    input n5047;
    input n5046;
    output \REG.mem_8_5 ;
    input n5045;
    input n5044;
    input n5043;
    input n5042;
    input n5041;
    input n5040;
    input n5039;
    input n5038;
    input n5037;
    input n5036;
    input n5035;
    output \REG.mem_7_10 ;
    input n5034;
    input n5033;
    input n5032;
    output \REG.mem_7_7 ;
    input n5031;
    input n5030;
    output \REG.mem_7_5 ;
    input n5029;
    input n5028;
    input n5027;
    input n5026;
    input n5025;
    output \REG.mem_7_0 ;
    input n5024;
    input n5023;
    input n5022;
    input n5021;
    input n5020;
    input n5019;
    output \REG.mem_6_10 ;
    input n5018;
    input n5017;
    input n5016;
    output \REG.mem_6_7 ;
    input n5015;
    input n5014;
    output \REG.mem_6_5 ;
    input n5013;
    input n5012;
    input n5011;
    input n5010;
    input n5009;
    output \REG.mem_6_0 ;
    input n5008;
    input n5007;
    input n5006;
    input n5005;
    input n5004;
    input n5003;
    output \REG.mem_5_10 ;
    input n5002;
    input n5001;
    input n5000;
    output \REG.mem_5_7 ;
    input n4999;
    input n4998;
    output \REG.mem_5_5 ;
    input n4997;
    input n4996;
    input n4995;
    input n4994;
    input n4993;
    output \REG.mem_5_0 ;
    input n4992;
    input n4991;
    input n4990;
    input n4989;
    input n4988;
    input n4987;
    output \REG.mem_4_10 ;
    input n4986;
    input n4985;
    input n4984;
    output \REG.mem_4_7 ;
    input n4983;
    input n4982;
    output \REG.mem_4_5 ;
    input n4981;
    input n4980;
    input n4979;
    input n4978;
    input n4977;
    output \REG.mem_4_0 ;
    input n4976;
    input n4975;
    input n4974;
    input n4973;
    input n4972;
    input n4971;
    output \REG.mem_3_10 ;
    input n4970;
    input n4969;
    output \REG.mem_3_8 ;
    output FT_OE_N_420;
    output n49;
    output n17;
    output n42;
    output n10;
    input n4968;
    output \REG.mem_3_7 ;
    input n4967;
    input n4966;
    output \REG.mem_3_5 ;
    input n4965;
    output n34;
    input n4964;
    input n4963;
    output n2;
    input n4962;
    input n4961;
    output \REG.mem_3_0 ;
    output n59;
    output n27;
    output n60;
    output n28;
    output n61;
    output n29;
    
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1 lscc_fifo_dc_inst (.rd_addr_r({Open_0, 
            Open_1, Open_2, Open_3, Open_4, Open_5, \rd_addr_r[0] }), 
            .\REG.mem_14_5 (\REG.mem_14_5 ), .\REG.mem_15_5 (\REG.mem_15_5 ), 
            .\dc32_fifo_data_in[6] (\dc32_fifo_data_in[6] ), .dc32_fifo_almost_full(dc32_fifo_almost_full), 
            .FIFO_CLK_c(FIFO_CLK_c), .reset_per_frame(reset_per_frame), 
            .\REG.mem_13_5 (\REG.mem_13_5 ), .\REG.mem_12_5 (\REG.mem_12_5 ), 
            .\dc32_fifo_data_in[5] (\dc32_fifo_data_in[5] ), .\dc32_fifo_data_in[4] (\dc32_fifo_data_in[4] ), 
            .\REG.mem_31_0 (\REG.mem_31_0 ), .GND_net(GND_net), .\dc32_fifo_data_in[3] (\dc32_fifo_data_in[3] ), 
            .\REG.mem_55_13 (\REG.mem_55_13 ), .\dc32_fifo_data_in[2] (\dc32_fifo_data_in[2] ), 
            .\REG.mem_38_7 (\REG.mem_38_7 ), .\REG.mem_39_7 (\REG.mem_39_7 ), 
            .\REG.mem_36_7 (\REG.mem_36_7 ), .\REG.mem_37_7 (\REG.mem_37_7 ), 
            .\REG.mem_16_8 (\REG.mem_16_8 ), .\REG.mem_18_8 (\REG.mem_18_8 ), 
            .\REG.mem_3_13 (\REG.mem_3_13 ), .\REG.mem_57_6 (\REG.mem_57_6 ), 
            .\dc32_fifo_data_in[1] (\dc32_fifo_data_in[1] ), .\REG.mem_63_11 (\REG.mem_63_11 ), 
            .\dc32_fifo_data_in[0] (\dc32_fifo_data_in[0] ), .\REG.mem_35_0 (\REG.mem_35_0 ), 
            .t_rd_fifo_en_w(t_rd_fifo_en_w), .\REG.out_raw[0] (\REG.out_raw[0] ), 
            .SLM_CLK_c(SLM_CLK_c), .\REG.mem_55_10 (\REG.mem_55_10 ), .n62(n62), 
            .n30(n30), .\REG.mem_31_3 (\REG.mem_31_3 ), .\REG.mem_48_7 (\REG.mem_48_7 ), 
            .\REG.mem_50_7 (\REG.mem_50_7 ), .\REG.mem_55_7 (\REG.mem_55_7 ), 
            .\REG.mem_48_10 (\REG.mem_48_10 ), .\REG.mem_50_10 (\REG.mem_50_10 ), 
            .wr_grey_sync_r({wr_grey_sync_r}), .\wr_addr_nxt_c[5] (\wr_addr_nxt_c[5] ), 
            .\REG.mem_23_8 (\REG.mem_23_8 ), .\REG.mem_25_5 (\REG.mem_25_5 ), 
            .\rd_grey_sync_r[0] (\rd_grey_sync_r[0] ), .\REG.mem_25_15 (\REG.mem_25_15 ), 
            .\REG.mem_14_12 (\REG.mem_14_12 ), .\REG.mem_15_12 (\REG.mem_15_12 ), 
            .DEBUG_3_c(DEBUG_3_c), .\REG.mem_13_12 (\REG.mem_13_12 ), .\REG.mem_12_12 (\REG.mem_12_12 ), 
            .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .dc32_fifo_almost_empty(dc32_fifo_almost_empty), .\REG.mem_6_1 (\REG.mem_6_1 ), 
            .\REG.mem_7_1 (\REG.mem_7_1 ), .\REG.mem_5_1 (\REG.mem_5_1 ), 
            .\REG.mem_4_1 (\REG.mem_4_1 ), .\REG.mem_57_9 (\REG.mem_57_9 ), 
            .\REG.mem_35_3 (\REG.mem_35_3 ), .\REG.mem_46_1 (\REG.mem_46_1 ), 
            .\REG.mem_47_1 (\REG.mem_47_1 ), .\REG.mem_45_1 (\REG.mem_45_1 ), 
            .\REG.mem_44_1 (\REG.mem_44_1 ), .\REG.mem_25_2 (\REG.mem_25_2 ), 
            .\dc32_fifo_data_in[15] (\dc32_fifo_data_in[15] ), .\dc32_fifo_data_in[14] (\dc32_fifo_data_in[14] ), 
            .\dc32_fifo_data_in[13] (\dc32_fifo_data_in[13] ), .\REG.mem_3_11 (\REG.mem_3_11 ), 
            .\REG.mem_31_2 (\REG.mem_31_2 ), .\REG.mem_50_12 (\REG.mem_50_12 ), 
            .\dc32_fifo_data_in[12] (\dc32_fifo_data_in[12] ), .\REG.mem_6_11 (\REG.mem_6_11 ), 
            .\REG.mem_7_11 (\REG.mem_7_11 ), .\REG.mem_5_11 (\REG.mem_5_11 ), 
            .\REG.mem_4_11 (\REG.mem_4_11 ), .\dc32_fifo_data_in[11] (\dc32_fifo_data_in[11] ), 
            .\REG.mem_48_12 (\REG.mem_48_12 ), .\REG.mem_3_4 (\REG.mem_3_4 ), 
            .\REG.mem_14_8 (\REG.mem_14_8 ), .\REG.mem_15_8 (\REG.mem_15_8 ), 
            .\REG.mem_8_14 (\REG.mem_8_14 ), .\REG.mem_9_14 (\REG.mem_9_14 ), 
            .\dc32_fifo_data_in[10] (\dc32_fifo_data_in[10] ), .\REG.mem_10_14 (\REG.mem_10_14 ), 
            .\REG.mem_11_14 (\REG.mem_11_14 ), .\REG.mem_63_6 (\REG.mem_63_6 ), 
            .\REG.mem_13_8 (\REG.mem_13_8 ), .\REG.mem_12_8 (\REG.mem_12_8 ), 
            .\REG.mem_14_14 (\REG.mem_14_14 ), .\REG.mem_15_14 (\REG.mem_15_14 ), 
            .\dc32_fifo_data_in[9] (\dc32_fifo_data_in[9] ), .\dc32_fifo_data_in[8] (\dc32_fifo_data_in[8] ), 
            .\REG.mem_3_1 (\REG.mem_3_1 ), .\dc32_fifo_data_in[7] (\dc32_fifo_data_in[7] ), 
            .\REG.mem_12_14 (\REG.mem_12_14 ), .\REG.mem_13_14 (\REG.mem_13_14 ), 
            .\REG.mem_42_8 (\REG.mem_42_8 ), .\REG.mem_43_8 (\REG.mem_43_8 ), 
            .\REG.mem_41_8 (\REG.mem_41_8 ), .\REG.mem_40_8 (\REG.mem_40_8 ), 
            .\REG.mem_18_12 (\REG.mem_18_12 ), .\REG.mem_16_12 (\REG.mem_16_12 ), 
            .\REG.mem_31_15 (\REG.mem_31_15 ), .\REG.mem_38_3 (\REG.mem_38_3 ), 
            .\REG.mem_39_3 (\REG.mem_39_3 ), .\REG.mem_37_3 (\REG.mem_37_3 ), 
            .\REG.mem_36_3 (\REG.mem_36_3 ), .\REG.mem_42_3 (\REG.mem_42_3 ), 
            .\REG.mem_43_3 (\REG.mem_43_3 ), .\REG.mem_14_7 (\REG.mem_14_7 ), 
            .\REG.mem_15_7 (\REG.mem_15_7 ), .\REG.mem_13_7 (\REG.mem_13_7 ), 
            .\REG.mem_12_7 (\REG.mem_12_7 ), .\REG.mem_41_3 (\REG.mem_41_3 ), 
            .\REG.mem_40_3 (\REG.mem_40_3 ), .\REG.mem_57_0 (\REG.mem_57_0 ), 
            .\REG.mem_10_11 (\REG.mem_10_11 ), .\REG.mem_11_11 (\REG.mem_11_11 ), 
            .\REG.mem_9_11 (\REG.mem_9_11 ), .\REG.mem_8_11 (\REG.mem_8_11 ), 
            .\REG.mem_63_12 (\REG.mem_63_12 ), .\REG.mem_55_12 (\REG.mem_55_12 ), 
            .\REG.mem_35_15 (\REG.mem_35_15 ), .\REG.mem_3_15 (\REG.mem_3_15 ), 
            .\wr_addr_nxt_c[3] (\wr_addr_nxt_c[3] ), .\REG.mem_50_9 (\REG.mem_50_9 ), 
            .\REG.mem_48_9 (\REG.mem_48_9 ), .\REG.mem_46_8 (\REG.mem_46_8 ), 
            .\REG.mem_47_8 (\REG.mem_47_8 ), .\REG.mem_46_3 (\REG.mem_46_3 ), 
            .\REG.mem_47_3 (\REG.mem_47_3 ), .\REG.mem_45_8 (\REG.mem_45_8 ), 
            .\REG.mem_44_8 (\REG.mem_44_8 ), .\REG.mem_16_2 (\REG.mem_16_2 ), 
            .\REG.mem_10_9 (\REG.mem_10_9 ), .\REG.mem_11_9 (\REG.mem_11_9 ), 
            .\REG.mem_45_3 (\REG.mem_45_3 ), .\REG.mem_44_3 (\REG.mem_44_3 ), 
            .\REG.mem_25_7 (\REG.mem_25_7 ), .\REG.mem_23_12 (\REG.mem_23_12 ), 
            .\REG.mem_18_2 (\REG.mem_18_2 ), .\REG.mem_38_0 (\REG.mem_38_0 ), 
            .\REG.mem_39_0 (\REG.mem_39_0 ), .\REG.mem_31_13 (\REG.mem_31_13 ), 
            .\REG.mem_37_0 (\REG.mem_37_0 ), .\REG.mem_36_0 (\REG.mem_36_0 ), 
            .\REG.mem_18_6 (\REG.mem_18_6 ), .\REG.mem_16_6 (\REG.mem_16_6 ), 
            .\REG.mem_9_9 (\REG.mem_9_9 ), .\REG.mem_8_9 (\REG.mem_8_9 ), 
            .\REG.mem_50_3 (\REG.mem_50_3 ), .\REG.mem_48_3 (\REG.mem_48_3 ), 
            .\REG.mem_42_0 (\REG.mem_42_0 ), .\REG.mem_43_0 (\REG.mem_43_0 ), 
            .\REG.mem_41_0 (\REG.mem_41_0 ), .\REG.mem_40_0 (\REG.mem_40_0 ), 
            .\REG.mem_14_11 (\REG.mem_14_11 ), .\REG.mem_15_11 (\REG.mem_15_11 ), 
            .\REG.mem_13_11 (\REG.mem_13_11 ), .\REG.mem_12_11 (\REG.mem_12_11 ), 
            .\REG.mem_38_5 (\REG.mem_38_5 ), .\REG.mem_39_5 (\REG.mem_39_5 ), 
            .\REG.mem_37_5 (\REG.mem_37_5 ), .\REG.mem_36_5 (\REG.mem_36_5 ), 
            .\REG.mem_57_13 (\REG.mem_57_13 ), .n6121(n6121), .VCC_net(VCC_net), 
            .\fifo_data_out[2] (\fifo_data_out[2] ), .n6118(n6118), .\fifo_data_out[1] (\fifo_data_out[1] ), 
            .\REG.mem_50_1 (\REG.mem_50_1 ), .\REG.mem_6_9 (\REG.mem_6_9 ), 
            .\REG.mem_7_9 (\REG.mem_7_9 ), .\REG.mem_48_1 (\REG.mem_48_1 ), 
            .n10556(n10556), .\fifo_data_out[3] (\fifo_data_out[3] ), .n10562(n10562), 
            .\fifo_data_out[4] (\fifo_data_out[4] ), .\REG.mem_18_11 (\REG.mem_18_11 ), 
            .\REG.mem_16_11 (\REG.mem_16_11 ), .\REG.mem_5_9 (\REG.mem_5_9 ), 
            .\REG.mem_4_9 (\REG.mem_4_9 ), .n10564(n10564), .\fifo_data_out[5] (\fifo_data_out[5] ), 
            .n10566(n10566), .\fifo_data_out[6] (\fifo_data_out[6] ), .n10568(n10568), 
            .\fifo_data_out[7] (\fifo_data_out[7] ), .n10570(n10570), .\fifo_data_out[8] (\fifo_data_out[8] ), 
            .n10572(n10572), .\fifo_data_out[9] (\fifo_data_out[9] ), .n10574(n10574), 
            .\fifo_data_out[10] (\fifo_data_out[10] ), .n10576(n10576), 
            .\fifo_data_out[11] (\fifo_data_out[11] ), .\REG.mem_31_5 (\REG.mem_31_5 ), 
            .n6085(n6085), .\fifo_data_out[0] (\fifo_data_out[0] ), .\REG.mem_25_12 (\REG.mem_25_12 ), 
            .\REG.mem_38_13 (\REG.mem_38_13 ), .\REG.mem_39_13 (\REG.mem_39_13 ), 
            .n10578(n10578), .\fifo_data_out[12] (\fifo_data_out[12] ), 
            .n10580(n10580), .\fifo_data_out[13] (\fifo_data_out[13] ), 
            .\rd_addr_r[6] (\rd_addr_r[6] ), .\REG.mem_6_15 (\REG.mem_6_15 ), 
            .\REG.mem_7_15 (\REG.mem_7_15 ), .n6045(n6045), .n6043(n6043), 
            .\REG.mem_5_15 (\REG.mem_5_15 ), .\REG.mem_4_15 (\REG.mem_4_15 ), 
            .\REG.mem_35_13 (\REG.mem_35_13 ), .n6024(n6024), .n6021(n6021), 
            .\REG.mem_63_15 (\REG.mem_63_15 ), .n6020(n6020), .\REG.mem_63_14 (\REG.mem_63_14 ), 
            .n6019(n6019), .\REG.mem_63_13 (\REG.mem_63_13 ), .n6018(n6018), 
            .n6017(n6017), .n6016(n6016), .\REG.mem_63_10 (\REG.mem_63_10 ), 
            .n6015(n6015), .\REG.mem_63_9 (\REG.mem_63_9 ), .n6014(n6014), 
            .\REG.mem_63_8 (\REG.mem_63_8 ), .n6013(n6013), .\REG.mem_63_7 (\REG.mem_63_7 ), 
            .n6012(n6012), .n6011(n6011), .\REG.mem_63_5 (\REG.mem_63_5 ), 
            .n6010(n6010), .\REG.mem_63_4 (\REG.mem_63_4 ), .n6009(n6009), 
            .\REG.mem_63_3 (\REG.mem_63_3 ), .n6008(n6008), .\REG.mem_63_2 (\REG.mem_63_2 ), 
            .n6007(n6007), .\REG.mem_63_1 (\REG.mem_63_1 ), .n6006(n6006), 
            .\REG.mem_63_0 (\REG.mem_63_0 ), .\REG.mem_25_6 (\REG.mem_25_6 ), 
            .\REG.mem_37_13 (\REG.mem_37_13 ), .\REG.mem_36_13 (\REG.mem_36_13 ), 
            .\REG.mem_57_4 (\REG.mem_57_4 ), .\REG.mem_18_7 (\REG.mem_18_7 ), 
            .\REG.mem_16_7 (\REG.mem_16_7 ), .\REG.mem_38_15 (\REG.mem_38_15 ), 
            .\REG.mem_39_15 (\REG.mem_39_15 ), .\REG.mem_23_11 (\REG.mem_23_11 ), 
            .\REG.mem_37_15 (\REG.mem_37_15 ), .\REG.mem_36_15 (\REG.mem_36_15 ), 
            .\REG.mem_25_11 (\REG.mem_25_11 ), .\REG.mem_57_12 (\REG.mem_57_12 ), 
            .\REG.mem_40_14 (\REG.mem_40_14 ), .\REG.mem_41_14 (\REG.mem_41_14 ), 
            .n5953(n5953), .rp_sync1_r({rp_sync1_r}), .\REG.mem_42_14 (\REG.mem_42_14 ), 
            .\REG.mem_43_14 (\REG.mem_43_14 ), .\REG.mem_46_14 (\REG.mem_46_14 ), 
            .\REG.mem_47_14 (\REG.mem_47_14 ), .n5952(n5952), .n5951(n5951), 
            .n5950(n5950), .n5949(n5949), .n5948(n5948), .n5947(n5947), 
            .n5946(n5946), .n5945(n5945), .\REG.mem_55_9 (\REG.mem_55_9 ), 
            .\REG.mem_44_14 (\REG.mem_44_14 ), .\REG.mem_45_14 (\REG.mem_45_14 ), 
            .\REG.mem_10_7 (\REG.mem_10_7 ), .\REG.mem_11_7 (\REG.mem_11_7 ), 
            .n5928(n5928), .n5927(n5927), .n5926(n5926), .n5924(n5924), 
            .n5923(n5923), .n5921(n5921), .\REG.mem_9_7 (\REG.mem_9_7 ), 
            .\REG.mem_8_7 (\REG.mem_8_7 ), .\REG.mem_40_4 (\REG.mem_40_4 ), 
            .\REG.mem_41_4 (\REG.mem_41_4 ), .\REG.mem_42_4 (\REG.mem_42_4 ), 
            .\REG.mem_43_4 (\REG.mem_43_4 ), .\REG.mem_46_4 (\REG.mem_46_4 ), 
            .\REG.mem_47_4 (\REG.mem_47_4 ), .\REG.mem_44_4 (\REG.mem_44_4 ), 
            .\REG.mem_45_4 (\REG.mem_45_4 ), .n5901(n5901), .\REG.mem_57_15 (\REG.mem_57_15 ), 
            .n5900(n5900), .\REG.mem_57_14 (\REG.mem_57_14 ), .n5899(n5899), 
            .n5898(n5898), .n5897(n5897), .\REG.mem_57_11 (\REG.mem_57_11 ), 
            .n5896(n5896), .\REG.mem_57_10 (\REG.mem_57_10 ), .n5895(n5895), 
            .n5894(n5894), .\REG.mem_57_8 (\REG.mem_57_8 ), .n5893(n5893), 
            .\REG.mem_57_7 (\REG.mem_57_7 ), .n5892(n5892), .n5891(n5891), 
            .\REG.mem_57_5 (\REG.mem_57_5 ), .n5890(n5890), .n5889(n5889), 
            .\REG.mem_57_3 (\REG.mem_57_3 ), .n5888(n5888), .\REG.mem_57_2 (\REG.mem_57_2 ), 
            .n5887(n5887), .\REG.mem_57_1 (\REG.mem_57_1 ), .\REG.mem_18_1 (\REG.mem_18_1 ), 
            .\REG.mem_16_1 (\REG.mem_16_1 ), .n5885(n5885), .\REG.mem_35_8 (\REG.mem_35_8 ), 
            .\REG.mem_38_8 (\REG.mem_38_8 ), .\REG.mem_39_8 (\REG.mem_39_8 ), 
            .\REG.mem_36_8 (\REG.mem_36_8 ), .\REG.mem_37_8 (\REG.mem_37_8 ), 
            .n5864(n5864), .wp_sync1_r({wp_sync1_r}), .n5863(n5863), .n5862(n5862), 
            .n5861(n5861), .n5860(n5860), .n5859(n5859), .n5858(n5858), 
            .\REG.mem_55_15 (\REG.mem_55_15 ), .n5857(n5857), .\REG.mem_55_14 (\REG.mem_55_14 ), 
            .n5856(n5856), .n5855(n5855), .n5854(n5854), .\REG.mem_55_11 (\REG.mem_55_11 ), 
            .n5853(n5853), .\rd_sig_diff0_w[0] (\rd_sig_diff0_w[0] ), .n5852(n5852), 
            .n5851(n5851), .\REG.mem_55_8 (\REG.mem_55_8 ), .n5850(n5850), 
            .n5849(n5849), .\REG.mem_55_6 (\REG.mem_55_6 ), .n5848(n5848), 
            .\REG.mem_55_5 (\REG.mem_55_5 ), .n5847(n5847), .\REG.mem_55_4 (\REG.mem_55_4 ), 
            .n5846(n5846), .\REG.mem_55_3 (\REG.mem_55_3 ), .n5845(n5845), 
            .\REG.mem_55_2 (\REG.mem_55_2 ), .n5844(n5844), .\REG.mem_55_1 (\REG.mem_55_1 ), 
            .n5843(n5843), .\REG.mem_55_0 (\REG.mem_55_0 ), .n5842(n5842), 
            .n5841(n5841), .n5839(n5839), .n5838(n5838), .n5837(n5837), 
            .\REG.mem_16_15 (\REG.mem_16_15 ), .\REG.mem_18_15 (\REG.mem_18_15 ), 
            .\REG.mem_23_15 (\REG.mem_23_15 ), .n5836(n5836), .\REG.mem_25_4 (\REG.mem_25_4 ), 
            .\REG.mem_35_2 (\REG.mem_35_2 ), .\REG.mem_31_4 (\REG.mem_31_4 ), 
            .\REG.mem_38_2 (\REG.mem_38_2 ), .\REG.mem_39_2 (\REG.mem_39_2 ), 
            .\REG.mem_36_2 (\REG.mem_36_2 ), .\REG.mem_37_2 (\REG.mem_37_2 ), 
            .\REG.mem_10_15 (\REG.mem_10_15 ), .\REG.mem_11_15 (\REG.mem_11_15 ), 
            .\REG.mem_48_2 (\REG.mem_48_2 ), .\REG.mem_50_2 (\REG.mem_50_2 ), 
            .\REG.mem_8_4 (\REG.mem_8_4 ), .\REG.mem_9_4 (\REG.mem_9_4 ), 
            .\REG.mem_10_4 (\REG.mem_10_4 ), .\REG.mem_11_4 (\REG.mem_11_4 ), 
            .n5771(n5771), .\REG.mem_50_15 (\REG.mem_50_15 ), .n5770(n5770), 
            .\REG.mem_50_14 (\REG.mem_50_14 ), .n5769(n5769), .\REG.mem_50_13 (\REG.mem_50_13 ), 
            .n5768(n5768), .n5767(n5767), .\REG.mem_50_11 (\REG.mem_50_11 ), 
            .n5766(n5766), .n5765(n5765), .n5764(n5764), .\REG.mem_50_8 (\REG.mem_50_8 ), 
            .n5763(n5763), .n5762(n5762), .\REG.mem_50_6 (\REG.mem_50_6 ), 
            .n5761(n5761), .\REG.mem_50_5 (\REG.mem_50_5 ), .n5760(n5760), 
            .\REG.mem_50_4 (\REG.mem_50_4 ), .n5759(n5759), .n5758(n5758), 
            .n5757(n5757), .\REG.mem_14_4 (\REG.mem_14_4 ), .\REG.mem_15_4 (\REG.mem_15_4 ), 
            .n10873(n10873), .\REG.mem_12_4 (\REG.mem_12_4 ), .\REG.mem_13_4 (\REG.mem_13_4 ), 
            .n10582(n10582), .\fifo_data_out[14] (\fifo_data_out[14] ), 
            .n10588(n10588), .\fifo_data_out[15] (\fifo_data_out[15] ), 
            .n5753(n5753), .\REG.mem_50_0 (\REG.mem_50_0 ), .\REG.mem_3_14 (\REG.mem_3_14 ), 
            .\REG.mem_6_14 (\REG.mem_6_14 ), .\REG.mem_7_14 (\REG.mem_7_14 ), 
            .\REG.mem_4_14 (\REG.mem_4_14 ), .\REG.mem_5_14 (\REG.mem_5_14 ), 
            .n5736(n5736), .\REG.mem_48_15 (\REG.mem_48_15 ), .n5735(n5735), 
            .\REG.mem_48_14 (\REG.mem_48_14 ), .n5734(n5734), .\REG.mem_48_13 (\REG.mem_48_13 ), 
            .n5733(n5733), .n5732(n5732), .\REG.mem_48_11 (\REG.mem_48_11 ), 
            .n5731(n5731), .n5730(n5730), .n5729(n5729), .\REG.mem_48_8 (\REG.mem_48_8 ), 
            .n5728(n5728), .n5727(n5727), .\REG.mem_48_6 (\REG.mem_48_6 ), 
            .n5726(n5726), .\REG.mem_48_5 (\REG.mem_48_5 ), .n5725(n5725), 
            .\REG.mem_48_4 (\REG.mem_48_4 ), .n5724(n5724), .n10877(n10877), 
            .\REG.mem_9_15 (\REG.mem_9_15 ), .\REG.mem_8_15 (\REG.mem_8_15 ), 
            .\REG.mem_31_7 (\REG.mem_31_7 ), .n5723(n5723), .n5722(n5722), 
            .n5721(n5721), .\REG.mem_48_0 (\REG.mem_48_0 ), .n5720(n5720), 
            .\REG.mem_47_15 (\REG.mem_47_15 ), .n5719(n5719), .n5718(n5718), 
            .\REG.mem_47_13 (\REG.mem_47_13 ), .n5717(n5717), .\REG.mem_47_12 (\REG.mem_47_12 ), 
            .n5716(n5716), .\REG.mem_47_11 (\REG.mem_47_11 ), .n5715(n5715), 
            .\REG.mem_47_10 (\REG.mem_47_10 ), .n5714(n5714), .\REG.mem_47_9 (\REG.mem_47_9 ), 
            .n5713(n5713), .n5712(n5712), .\REG.mem_47_7 (\REG.mem_47_7 ), 
            .n5711(n5711), .\REG.mem_47_6 (\REG.mem_47_6 ), .n5710(n5710), 
            .\REG.mem_47_5 (\REG.mem_47_5 ), .n5709(n5709), .n5708(n5708), 
            .n5707(n5707), .\REG.mem_47_2 (\REG.mem_47_2 ), .n5706(n5706), 
            .n5705(n5705), .\REG.mem_47_0 (\REG.mem_47_0 ), .n5704(n5704), 
            .\REG.mem_46_15 (\REG.mem_46_15 ), .n5703(n5703), .\REG.mem_31_12 (\REG.mem_31_12 ), 
            .n5702(n5702), .\REG.mem_46_13 (\REG.mem_46_13 ), .n5701(n5701), 
            .\REG.mem_46_12 (\REG.mem_46_12 ), .n5700(n5700), .\REG.mem_46_11 (\REG.mem_46_11 ), 
            .n5699(n5699), .\REG.mem_46_10 (\REG.mem_46_10 ), .n5698(n5698), 
            .\REG.mem_46_9 (\REG.mem_46_9 ), .n5697(n5697), .n5696(n5696), 
            .\REG.mem_46_7 (\REG.mem_46_7 ), .n5695(n5695), .\REG.mem_46_6 (\REG.mem_46_6 ), 
            .n5694(n5694), .\REG.mem_46_5 (\REG.mem_46_5 ), .n5693(n5693), 
            .n5692(n5692), .n5691(n5691), .\REG.mem_46_2 (\REG.mem_46_2 ), 
            .n5690(n5690), .n5689(n5689), .\REG.mem_46_0 (\REG.mem_46_0 ), 
            .n5688(n5688), .\REG.mem_45_15 (\REG.mem_45_15 ), .n5687(n5687), 
            .n5686(n5686), .\REG.mem_45_13 (\REG.mem_45_13 ), .n5685(n5685), 
            .\REG.mem_45_12 (\REG.mem_45_12 ), .n5684(n5684), .\REG.mem_45_11 (\REG.mem_45_11 ), 
            .n5683(n5683), .\REG.mem_45_10 (\REG.mem_45_10 ), .n5682(n5682), 
            .\REG.mem_45_9 (\REG.mem_45_9 ), .n5681(n5681), .n5680(n5680), 
            .\REG.mem_45_7 (\REG.mem_45_7 ), .n5679(n5679), .\REG.mem_45_6 (\REG.mem_45_6 ), 
            .n5678(n5678), .\REG.mem_45_5 (\REG.mem_45_5 ), .\REG.mem_38_6 (\REG.mem_38_6 ), 
            .\REG.mem_39_6 (\REG.mem_39_6 ), .\REG.mem_37_6 (\REG.mem_37_6 ), 
            .\REG.mem_36_6 (\REG.mem_36_6 ), .n5677(n5677), .\REG.mem_31_11 (\REG.mem_31_11 ), 
            .n5676(n5676), .\REG.mem_42_5 (\REG.mem_42_5 ), .\REG.mem_43_5 (\REG.mem_43_5 ), 
            .n5675(n5675), .\REG.mem_45_2 (\REG.mem_45_2 ), .n5674(n5674), 
            .n5673(n5673), .\REG.mem_45_0 (\REG.mem_45_0 ), .n5671(n5671), 
            .\REG.mem_44_15 (\REG.mem_44_15 ), .n5670(n5670), .n5669(n5669), 
            .\REG.mem_44_13 (\REG.mem_44_13 ), .n5668(n5668), .\REG.mem_44_12 (\REG.mem_44_12 ), 
            .n5666(n5666), .\REG.mem_44_11 (\REG.mem_44_11 ), .n5665(n5665), 
            .\REG.mem_44_10 (\REG.mem_44_10 ), .n5664(n5664), .\REG.mem_44_9 (\REG.mem_44_9 ), 
            .n5662(n5662), .n5661(n5661), .\REG.mem_44_7 (\REG.mem_44_7 ), 
            .n5660(n5660), .\REG.mem_44_6 (\REG.mem_44_6 ), .n5659(n5659), 
            .\REG.mem_44_5 (\REG.mem_44_5 ), .n5658(n5658), .n5657(n5657), 
            .n5656(n5656), .\REG.mem_44_2 (\REG.mem_44_2 ), .n5655(n5655), 
            .n5654(n5654), .\REG.mem_44_0 (\REG.mem_44_0 ), .n5653(n5653), 
            .\REG.mem_43_15 (\REG.mem_43_15 ), .n5652(n5652), .n5651(n5651), 
            .\REG.mem_43_13 (\REG.mem_43_13 ), .n5650(n5650), .\REG.mem_43_12 (\REG.mem_43_12 ), 
            .n5649(n5649), .\REG.mem_43_11 (\REG.mem_43_11 ), .n5648(n5648), 
            .\REG.mem_43_10 (\REG.mem_43_10 ), .n5647(n5647), .\REG.mem_43_9 (\REG.mem_43_9 ), 
            .n5646(n5646), .n5645(n5645), .\REG.mem_43_7 (\REG.mem_43_7 ), 
            .n5644(n5644), .\REG.mem_43_6 (\REG.mem_43_6 ), .\REG.mem_41_5 (\REG.mem_41_5 ), 
            .\REG.mem_40_5 (\REG.mem_40_5 ), .\REG.mem_23_1 (\REG.mem_23_1 ), 
            .\rd_addr_p1_w[0] (\rd_addr_p1_w[0] ), .\REG.mem_35_11 (\REG.mem_35_11 ), 
            .n5643(n5643), .n5642(n5642), .n5641(n5641), .n5640(n5640), 
            .\REG.mem_43_2 (\REG.mem_43_2 ), .n5639(n5639), .\REG.mem_43_1 (\REG.mem_43_1 ), 
            .n5638(n5638), .n5637(n5637), .\REG.mem_42_15 (\REG.mem_42_15 ), 
            .n5636(n5636), .n5635(n5635), .\REG.mem_42_13 (\REG.mem_42_13 ), 
            .n5634(n5634), .\REG.mem_42_12 (\REG.mem_42_12 ), .n5633(n5633), 
            .\REG.mem_42_11 (\REG.mem_42_11 ), .n5632(n5632), .\REG.mem_42_10 (\REG.mem_42_10 ), 
            .n5631(n5631), .\REG.mem_42_9 (\REG.mem_42_9 ), .n5630(n5630), 
            .n5629(n5629), .\REG.mem_42_7 (\REG.mem_42_7 ), .n4916(n4916), 
            .\REG.mem_31_6 (\REG.mem_31_6 ), .\REG.mem_23_2 (\REG.mem_23_2 ), 
            .\REG.mem_38_11 (\REG.mem_38_11 ), .\REG.mem_39_11 (\REG.mem_39_11 ), 
            .\REG.mem_37_11 (\REG.mem_37_11 ), .\REG.mem_36_11 (\REG.mem_36_11 ), 
            .n5628(n5628), .\REG.mem_42_6 (\REG.mem_42_6 ), .n5627(n5627), 
            .n5626(n5626), .n5625(n5625), .n5624(n5624), .\REG.mem_42_2 (\REG.mem_42_2 ), 
            .n5623(n5623), .\REG.mem_42_1 (\REG.mem_42_1 ), .n5622(n5622), 
            .n5621(n5621), .\REG.mem_41_15 (\REG.mem_41_15 ), .n5620(n5620), 
            .n5619(n5619), .\REG.mem_41_13 (\REG.mem_41_13 ), .n5618(n5618), 
            .\REG.mem_41_12 (\REG.mem_41_12 ), .n5617(n5617), .\REG.mem_41_11 (\REG.mem_41_11 ), 
            .n5616(n5616), .\REG.mem_41_10 (\REG.mem_41_10 ), .n5615(n5615), 
            .\REG.mem_41_9 (\REG.mem_41_9 ), .n5614(n5614), .n5613(n5613), 
            .\REG.mem_41_7 (\REG.mem_41_7 ), .\REG.mem_3_2 (\REG.mem_3_2 ), 
            .n5612(n5612), .\REG.mem_41_6 (\REG.mem_41_6 ), .n5611(n5611), 
            .n5610(n5610), .n5609(n5609), .n5608(n5608), .\REG.mem_41_2 (\REG.mem_41_2 ), 
            .n5607(n5607), .\REG.mem_41_1 (\REG.mem_41_1 ), .n5606(n5606), 
            .n5605(n5605), .\REG.mem_40_15 (\REG.mem_40_15 ), .n5604(n5604), 
            .n5603(n5603), .\REG.mem_40_13 (\REG.mem_40_13 ), .n5602(n5602), 
            .\REG.mem_40_12 (\REG.mem_40_12 ), .n5601(n5601), .\REG.mem_40_11 (\REG.mem_40_11 ), 
            .n5600(n5600), .\REG.mem_40_10 (\REG.mem_40_10 ), .n5599(n5599), 
            .\REG.mem_40_9 (\REG.mem_40_9 ), .n5598(n5598), .n5597(n5597), 
            .\REG.mem_40_7 (\REG.mem_40_7 ), .\REG.mem_25_9 (\REG.mem_25_9 ), 
            .n4904(n4904), .n4903(n4903), .n4901(n4901), .n4899(n4899), 
            .n5596(n5596), .\REG.mem_40_6 (\REG.mem_40_6 ), .n5595(n5595), 
            .n5594(n5594), .n5593(n5593), .n5592(n5592), .\REG.mem_40_2 (\REG.mem_40_2 ), 
            .n5591(n5591), .\REG.mem_40_1 (\REG.mem_40_1 ), .n5590(n5590), 
            .n5589(n5589), .n5588(n5588), .\REG.mem_39_14 (\REG.mem_39_14 ), 
            .n5587(n5587), .n5586(n5586), .\REG.mem_39_12 (\REG.mem_39_12 ), 
            .n5585(n5585), .n5584(n5584), .\REG.mem_39_10 (\REG.mem_39_10 ), 
            .n5583(n5583), .\REG.mem_39_9 (\REG.mem_39_9 ), .n5582(n5582), 
            .n5581(n5581), .n4898(n4898), .\REG.mem_14_1 (\REG.mem_14_1 ), 
            .\REG.mem_15_1 (\REG.mem_15_1 ), .DEBUG_5_c(DEBUG_5_c), .\REG.mem_13_1 (\REG.mem_13_1 ), 
            .\REG.mem_12_1 (\REG.mem_12_1 ), .\REG.mem_3_3 (\REG.mem_3_3 ), 
            .n5580(n5580), .n5579(n5579), .n5578(n5578), .\REG.mem_39_4 (\REG.mem_39_4 ), 
            .n5577(n5577), .n5576(n5576), .n5575(n5575), .\REG.mem_39_1 (\REG.mem_39_1 ), 
            .n5573(n5573), .n5572(n5572), .n5571(n5571), .\REG.mem_38_14 (\REG.mem_38_14 ), 
            .n5570(n5570), .n5569(n5569), .\REG.mem_38_12 (\REG.mem_38_12 ), 
            .n5568(n5568), .n5567(n5567), .\REG.mem_38_10 (\REG.mem_38_10 ), 
            .n5566(n5566), .\REG.mem_38_9 (\REG.mem_38_9 ), .n5565(n5565), 
            .n5564(n5564), .n5563(n5563), .n5562(n5562), .n5561(n5561), 
            .\REG.mem_38_4 (\REG.mem_38_4 ), .n5560(n5560), .n5559(n5559), 
            .n5558(n5558), .\REG.mem_38_1 (\REG.mem_38_1 ), .n5556(n5556), 
            .n5555(n5555), .n5554(n5554), .\REG.mem_37_14 (\REG.mem_37_14 ), 
            .n5553(n5553), .n5552(n5552), .\REG.mem_37_12 (\REG.mem_37_12 ), 
            .n5551(n5551), .n5550(n5550), .\REG.mem_37_10 (\REG.mem_37_10 ), 
            .n5549(n5549), .\REG.mem_37_9 (\REG.mem_37_9 ), .\REG.mem_25_13 (\REG.mem_25_13 ), 
            .\REG.out_raw[15] (\REG.out_raw[15] ), .\REG.out_raw[14] (\REG.out_raw[14] ), 
            .\REG.out_raw[13] (\REG.out_raw[13] ), .\REG.out_raw[12] (\REG.out_raw[12] ), 
            .\REG.out_raw[11] (\REG.out_raw[11] ), .n5548(n5548), .n5547(n5547), 
            .n5546(n5546), .n5545(n5545), .n5544(n5544), .\REG.mem_37_4 (\REG.mem_37_4 ), 
            .n5543(n5543), .n5542(n5542), .n5541(n5541), .\REG.mem_37_1 (\REG.mem_37_1 ), 
            .n5540(n5540), .\REG.out_raw[10] (\REG.out_raw[10] ), .\REG.out_raw[9] (\REG.out_raw[9] ), 
            .\REG.out_raw[8] (\REG.out_raw[8] ), .\REG.out_raw[7] (\REG.out_raw[7] ), 
            .\REG.out_raw[6] (\REG.out_raw[6] ), .\REG.out_raw[5] (\REG.out_raw[5] ), 
            .\REG.out_raw[4] (\REG.out_raw[4] ), .\REG.out_raw[3] (\REG.out_raw[3] ), 
            .\REG.out_raw[2] (\REG.out_raw[2] ), .\REG.out_raw[1] (\REG.out_raw[1] ), 
            .n5526(n5526), .n5525(n5525), .\REG.mem_36_14 (\REG.mem_36_14 ), 
            .n5524(n5524), .n5523(n5523), .\REG.mem_36_12 (\REG.mem_36_12 ), 
            .n5522(n5522), .n5521(n5521), .\REG.mem_36_10 (\REG.mem_36_10 ), 
            .n5520(n5520), .\REG.mem_36_9 (\REG.mem_36_9 ), .n5519(n5519), 
            .n5518(n5518), .n5517(n5517), .n5516(n5516), .\rd_sig_diff0_w[2] (\rd_sig_diff0_w[2] ), 
            .n5515(n5515), .\REG.mem_36_4 (\REG.mem_36_4 ), .n5514(n5514), 
            .n5513(n5513), .n5512(n5512), .\REG.mem_36_1 (\REG.mem_36_1 ), 
            .n5511(n5511), .n5507(n5507), .n5506(n5506), .\REG.mem_35_14 (\REG.mem_35_14 ), 
            .n5505(n5505), .n5504(n5504), .\REG.mem_35_12 (\REG.mem_35_12 ), 
            .n5503(n5503), .n5502(n5502), .\REG.mem_35_10 (\REG.mem_35_10 ), 
            .n5501(n5501), .\REG.mem_35_9 (\REG.mem_35_9 ), .n5500(n5500), 
            .\rd_sig_diff0_w[1] (\rd_sig_diff0_w[1] ), .n5499(n5499), .\REG.mem_35_7 (\REG.mem_35_7 ), 
            .n5498(n5498), .\REG.mem_35_6 (\REG.mem_35_6 ), .n5497(n5497), 
            .\REG.mem_35_5 (\REG.mem_35_5 ), .n5496(n5496), .\REG.mem_35_4 (\REG.mem_35_4 ), 
            .n5495(n5495), .n5494(n5494), .n5493(n5493), .\REG.mem_35_1 (\REG.mem_35_1 ), 
            .n5492(n5492), .\REG.mem_6_3 (\REG.mem_6_3 ), .\REG.mem_7_3 (\REG.mem_7_3 ), 
            .\REG.mem_5_3 (\REG.mem_5_3 ), .\REG.mem_4_3 (\REG.mem_4_3 ), 
            .n5441(n5441), .n5440(n5440), .\REG.mem_31_14 (\REG.mem_31_14 ), 
            .n5439(n5439), .n5438(n5438), .n5437(n5437), .\REG.mem_25_1 (\REG.mem_25_1 ), 
            .n5436(n5436), .\REG.mem_31_10 (\REG.mem_31_10 ), .n58(n58), 
            .n5435(n5435), .\REG.mem_31_9 (\REG.mem_31_9 ), .n5434(n5434), 
            .\REG.mem_31_8 (\REG.mem_31_8 ), .n5433(n5433), .n5432(n5432), 
            .n5431(n5431), .n5430(n5430), .n5429(n5429), .n5428(n5428), 
            .n5427(n5427), .\REG.mem_31_1 (\REG.mem_31_1 ), .n5426(n5426), 
            .n26(n26), .DEBUG_1_c_c(DEBUG_1_c_c), .write_to_dc32_fifo_latched_N_425(write_to_dc32_fifo_latched_N_425), 
            .n5345(n5345), .n5344(n5344), .\REG.mem_25_14 (\REG.mem_25_14 ), 
            .n5343(n5343), .n5342(n5342), .n5341(n5341), .n5340(n5340), 
            .\REG.mem_25_10 (\REG.mem_25_10 ), .n5339(n5339), .n5338(n5338), 
            .\REG.mem_25_8 (\REG.mem_25_8 ), .n5337(n5337), .n5336(n5336), 
            .n5335(n5335), .n5334(n5334), .n5333(n5333), .\REG.mem_25_3 (\REG.mem_25_3 ), 
            .n5332(n5332), .n5331(n5331), .n5330(n5330), .\REG.mem_25_0 (\REG.mem_25_0 ), 
            .\REG.mem_14_15 (\REG.mem_14_15 ), .\REG.mem_15_15 (\REG.mem_15_15 ), 
            .\REG.mem_6_13 (\REG.mem_6_13 ), .\REG.mem_7_13 (\REG.mem_7_13 ), 
            .n5306(n5306), .n5305(n5305), .\REG.mem_23_14 (\REG.mem_23_14 ), 
            .n5304(n5304), .\REG.mem_23_13 (\REG.mem_23_13 ), .n5303(n5303), 
            .n5302(n5302), .n5301(n5301), .\REG.mem_23_10 (\REG.mem_23_10 ), 
            .n5300(n5300), .\REG.mem_23_9 (\REG.mem_23_9 ), .n5299(n5299), 
            .n5298(n5298), .\REG.mem_23_7 (\REG.mem_23_7 ), .n5297(n5297), 
            .\REG.mem_23_6 (\REG.mem_23_6 ), .n5296(n5296), .\REG.mem_23_5 (\REG.mem_23_5 ), 
            .n5295(n5295), .\REG.mem_23_4 (\REG.mem_23_4 ), .n5294(n5294), 
            .\REG.mem_23_3 (\REG.mem_23_3 ), .n5293(n5293), .n5292(n5292), 
            .n5290(n5290), .\REG.mem_23_0 (\REG.mem_23_0 ), .\rd_grey_sync_r[5] (\rd_grey_sync_r[5] ), 
            .\REG.mem_5_13 (\REG.mem_5_13 ), .\REG.mem_4_13 (\REG.mem_4_13 ), 
            .\rd_grey_sync_r[4] (\rd_grey_sync_r[4] ), .\rd_grey_sync_r[3] (\rd_grey_sync_r[3] ), 
            .\rd_grey_sync_r[2] (\rd_grey_sync_r[2] ), .\rd_grey_sync_r[1] (\rd_grey_sync_r[1] ), 
            .\REG.mem_13_15 (\REG.mem_13_15 ), .\REG.mem_12_15 (\REG.mem_12_15 ), 
            .n51(n51), .n19(n19), .\wr_addr_nxt_c[1] (\wr_addr_nxt_c[1] ), 
            .\REG.mem_10_0 (\REG.mem_10_0 ), .\REG.mem_11_0 (\REG.mem_11_0 ), 
            .\REG.mem_10_3 (\REG.mem_10_3 ), .\REG.mem_11_3 (\REG.mem_11_3 ), 
            .n5224(n5224), .n5223(n5223), .\REG.mem_18_14 (\REG.mem_18_14 ), 
            .n5222(n5222), .\REG.mem_18_13 (\REG.mem_18_13 ), .n5221(n5221), 
            .n5220(n5220), .\REG.mem_9_3 (\REG.mem_9_3 ), .\REG.mem_8_3 (\REG.mem_8_3 ), 
            .\REG.mem_9_0 (\REG.mem_9_0 ), .\REG.mem_8_0 (\REG.mem_8_0 ), 
            .\REG.mem_10_13 (\REG.mem_10_13 ), .\REG.mem_11_13 (\REG.mem_11_13 ), 
            .n52(n52), .\REG.mem_9_13 (\REG.mem_9_13 ), .\REG.mem_8_13 (\REG.mem_8_13 ), 
            .n20(n20), .n5219(n5219), .\REG.mem_18_10 (\REG.mem_18_10 ), 
            .n5218(n5218), .\REG.mem_18_9 (\REG.mem_18_9 ), .n5217(n5217), 
            .n5216(n5216), .n5215(n5215), .n5214(n5214), .\REG.mem_18_5 (\REG.mem_18_5 ), 
            .n5213(n5213), .\REG.mem_18_4 (\REG.mem_18_4 ), .n5212(n5212), 
            .\REG.mem_18_3 (\REG.mem_18_3 ), .n5211(n5211), .n5210(n5210), 
            .n5209(n5209), .\REG.mem_18_0 (\REG.mem_18_0 ), .\REG.mem_14_13 (\REG.mem_14_13 ), 
            .\REG.mem_15_13 (\REG.mem_15_13 ), .\REG.mem_13_13 (\REG.mem_13_13 ), 
            .\REG.mem_12_13 (\REG.mem_12_13 ), .\REG.mem_6_4 (\REG.mem_6_4 ), 
            .\REG.mem_7_4 (\REG.mem_7_4 ), .\REG.mem_5_4 (\REG.mem_5_4 ), 
            .\REG.mem_4_4 (\REG.mem_4_4 ), .get_next_word(get_next_word), 
            .n5188(n5188), .n5186(n5186), .\REG.mem_16_14 (\REG.mem_16_14 ), 
            .n5185(n5185), .\REG.mem_16_13 (\REG.mem_16_13 ), .\REG.mem_6_8 (\REG.mem_6_8 ), 
            .\REG.mem_7_8 (\REG.mem_7_8 ), .\REG.mem_3_6 (\REG.mem_3_6 ), 
            .n5184(n5184), .\REG.mem_5_8 (\REG.mem_5_8 ), .\REG.mem_4_8 (\REG.mem_4_8 ), 
            .\REG.mem_6_2 (\REG.mem_6_2 ), .\REG.mem_7_2 (\REG.mem_7_2 ), 
            .\REG.mem_5_2 (\REG.mem_5_2 ), .\REG.mem_4_2 (\REG.mem_4_2 ), 
            .rd_fifo_en_w(rd_fifo_en_w), .n5183(n5183), .n5182(n5182), 
            .\REG.mem_16_10 (\REG.mem_16_10 ), .n5181(n5181), .\REG.mem_16_9 (\REG.mem_16_9 ), 
            .n5180(n5180), .n5179(n5179), .n5178(n5178), .n5177(n5177), 
            .\REG.mem_16_5 (\REG.mem_16_5 ), .n5176(n5176), .\REG.mem_16_4 (\REG.mem_16_4 ), 
            .\REG.mem_3_12 (\REG.mem_3_12 ), .n5175(n5175), .\REG.mem_16_3 (\REG.mem_16_3 ), 
            .n5174(n5174), .n5173(n5173), .n5172(n5172), .\REG.mem_16_0 (\REG.mem_16_0 ), 
            .n5169(n5169), .n5168(n5168), .n5167(n5167), .n47(n47), 
            .n5166(n5166), .n15(n15), .n5165(n5165), .n5164(n5164), 
            .\REG.mem_15_10 (\REG.mem_15_10 ), .n5163(n5163), .\REG.mem_15_9 (\REG.mem_15_9 ), 
            .n5162(n5162), .n5161(n5161), .n5160(n5160), .\REG.mem_15_6 (\REG.mem_15_6 ), 
            .n5159(n5159), .n5158(n5158), .n5157(n5157), .\REG.mem_15_3 (\REG.mem_15_3 ), 
            .n5156(n5156), .\REG.mem_15_2 (\REG.mem_15_2 ), .n5155(n5155), 
            .n5154(n5154), .\REG.mem_15_0 (\REG.mem_15_0 ), .n5153(n5153), 
            .n5152(n5152), .\REG.mem_6_6 (\REG.mem_6_6 ), .\REG.mem_7_6 (\REG.mem_7_6 ), 
            .n5151(n5151), .n5150(n5150), .n5149(n5149), .n5148(n5148), 
            .\REG.mem_14_10 (\REG.mem_14_10 ), .n5147(n5147), .\REG.mem_14_9 (\REG.mem_14_9 ), 
            .n5146(n5146), .n5145(n5145), .n5144(n5144), .\REG.mem_14_6 (\REG.mem_14_6 ), 
            .\REG.mem_4_6 (\REG.mem_4_6 ), .\REG.mem_5_6 (\REG.mem_5_6 ), 
            .n5143(n5143), .n5142(n5142), .n5141(n5141), .\REG.mem_14_3 (\REG.mem_14_3 ), 
            .n5140(n5140), .\REG.mem_14_2 (\REG.mem_14_2 ), .n5139(n5139), 
            .n5138(n5138), .\REG.mem_14_0 (\REG.mem_14_0 ), .n5137(n5137), 
            .n5136(n5136), .n5135(n5135), .n5134(n5134), .n5133(n5133), 
            .n5132(n5132), .\REG.mem_13_10 (\REG.mem_13_10 ), .\REG.mem_13_9 (\REG.mem_13_9 ), 
            .\REG.mem_12_9 (\REG.mem_12_9 ), .n5131(n5131), .n5130(n5130), 
            .n5129(n5129), .n5128(n5128), .\REG.mem_13_6 (\REG.mem_13_6 ), 
            .n5127(n5127), .n5126(n5126), .n5125(n5125), .\REG.mem_13_3 (\REG.mem_13_3 ), 
            .n5124(n5124), .\REG.mem_13_2 (\REG.mem_13_2 ), .n5123(n5123), 
            .\REG.mem_10_8 (\REG.mem_10_8 ), .\REG.mem_11_8 (\REG.mem_11_8 ), 
            .n5122(n5122), .\REG.mem_13_0 (\REG.mem_13_0 ), .n5121(n5121), 
            .n5120(n5120), .n5119(n5119), .n5118(n5118), .\REG.mem_3_9 (\REG.mem_3_9 ), 
            .\REG.mem_9_8 (\REG.mem_9_8 ), .\REG.mem_8_8 (\REG.mem_8_8 ), 
            .n5117(n5117), .\REG.mem_8_6 (\REG.mem_8_6 ), .\REG.mem_9_6 (\REG.mem_9_6 ), 
            .n5116(n5116), .\REG.mem_12_10 (\REG.mem_12_10 ), .\REG.mem_10_6 (\REG.mem_10_6 ), 
            .\REG.mem_11_6 (\REG.mem_11_6 ), .n53(n53), .n21(n21), .n5115(n5115), 
            .n5114(n5114), .n5113(n5113), .n5112(n5112), .\REG.mem_12_6 (\REG.mem_12_6 ), 
            .n50(n50), .n5111(n5111), .n18(n18), .\REG.mem_6_12 (\REG.mem_6_12 ), 
            .\REG.mem_7_12 (\REG.mem_7_12 ), .n5110(n5110), .n5109(n5109), 
            .\REG.mem_12_3 (\REG.mem_12_3 ), .n5108(n5108), .\REG.mem_12_2 (\REG.mem_12_2 ), 
            .\REG.mem_4_12 (\REG.mem_4_12 ), .\REG.mem_5_12 (\REG.mem_5_12 ), 
            .\REG.mem_10_2 (\REG.mem_10_2 ), .\REG.mem_11_2 (\REG.mem_11_2 ), 
            .n5107(n5107), .\REG.mem_9_2 (\REG.mem_9_2 ), .\REG.mem_8_2 (\REG.mem_8_2 ), 
            .n54(n54), .n22(n22), .n5106(n5106), .\REG.mem_12_0 (\REG.mem_12_0 ), 
            .\rd_addr_nxt_c_6__N_498[3] (\rd_addr_nxt_c_6__N_498[3] ), .n5105(n5105), 
            .n5104(n5104), .n5103(n5103), .n5102(n5102), .\REG.mem_11_12 (\REG.mem_11_12 ), 
            .n5101(n5101), .n5100(n5100), .\REG.mem_11_10 (\REG.mem_11_10 ), 
            .n5099(n5099), .n5098(n5098), .n5097(n5097), .n5096(n5096), 
            .n5095(n5095), .\REG.mem_11_5 (\REG.mem_11_5 ), .n5094(n5094), 
            .n5093(n5093), .n5092(n5092), .n5091(n5091), .\REG.mem_11_1 (\REG.mem_11_1 ), 
            .n5090(n5090), .n5089(n5089), .n5088(n5088), .\rd_addr_nxt_c_6__N_498[5] (\rd_addr_nxt_c_6__N_498[5] ), 
            .n5087(n5087), .n5086(n5086), .\REG.mem_10_12 (\REG.mem_10_12 ), 
            .n5085(n5085), .n5084(n5084), .\REG.mem_10_10 (\REG.mem_10_10 ), 
            .n5083(n5083), .n5082(n5082), .n5081(n5081), .n5080(n5080), 
            .n5079(n5079), .\REG.mem_10_5 (\REG.mem_10_5 ), .\REG.mem_10_1 (\REG.mem_10_1 ), 
            .\REG.mem_9_1 (\REG.mem_9_1 ), .\REG.mem_8_1 (\REG.mem_8_1 ), 
            .\rd_addr_nxt_c_6__N_498[2] (\rd_addr_nxt_c_6__N_498[2] ), .n56(n56), 
            .n24(n24), .n5078(n5078), .n55(n55), .n23(n23), .n5077(n5077), 
            .n40(n40), .n8(n8), .n5076(n5076), .n5075(n5075), .n5074(n5074), 
            .n5073(n5073), .n5072(n5072), .n5071(n5071), .n5070(n5070), 
            .\REG.mem_9_12 (\REG.mem_9_12 ), .n5069(n5069), .n5068(n5068), 
            .\REG.mem_9_10 (\REG.mem_9_10 ), .n5067(n5067), .n5066(n5066), 
            .n5065(n5065), .n57(n57), .n5064(n5064), .n25(n25), .n5063(n5063), 
            .\REG.mem_9_5 (\REG.mem_9_5 ), .n5062(n5062), .n5061(n5061), 
            .n5060(n5060), .n5059(n5059), .n5057(n5057), .n5056(n5056), 
            .n5055(n5055), .n5054(n5054), .n5053(n5053), .\REG.mem_8_12 (\REG.mem_8_12 ), 
            .n5052(n5052), .n5051(n5051), .\REG.mem_8_10 (\REG.mem_8_10 ), 
            .n5050(n5050), .n5049(n5049), .n5048(n5048), .n5047(n5047), 
            .n5046(n5046), .\REG.mem_8_5 (\REG.mem_8_5 ), .n5045(n5045), 
            .n5044(n5044), .n5043(n5043), .n5042(n5042), .n5041(n5041), 
            .n5040(n5040), .n5039(n5039), .n5038(n5038), .n5037(n5037), 
            .n5036(n5036), .n5035(n5035), .\REG.mem_7_10 (\REG.mem_7_10 ), 
            .n5034(n5034), .n5033(n5033), .n5032(n5032), .\REG.mem_7_7 (\REG.mem_7_7 ), 
            .n5031(n5031), .n5030(n5030), .\REG.mem_7_5 (\REG.mem_7_5 ), 
            .n5029(n5029), .n5028(n5028), .n5027(n5027), .n5026(n5026), 
            .n5025(n5025), .\REG.mem_7_0 (\REG.mem_7_0 ), .n5024(n5024), 
            .n5023(n5023), .n5022(n5022), .n5021(n5021), .n5020(n5020), 
            .n5019(n5019), .\REG.mem_6_10 (\REG.mem_6_10 ), .n5018(n5018), 
            .n5017(n5017), .n5016(n5016), .\REG.mem_6_7 (\REG.mem_6_7 ), 
            .n5015(n5015), .n5014(n5014), .\REG.mem_6_5 (\REG.mem_6_5 ), 
            .n5013(n5013), .n5012(n5012), .n5011(n5011), .n5010(n5010), 
            .n5009(n5009), .\REG.mem_6_0 (\REG.mem_6_0 ), .n5008(n5008), 
            .n5007(n5007), .n5006(n5006), .n5005(n5005), .n5004(n5004), 
            .n5003(n5003), .\REG.mem_5_10 (\REG.mem_5_10 ), .n5002(n5002), 
            .n5001(n5001), .n5000(n5000), .\REG.mem_5_7 (\REG.mem_5_7 ), 
            .n4999(n4999), .n4998(n4998), .\REG.mem_5_5 (\REG.mem_5_5 ), 
            .n4997(n4997), .n4996(n4996), .n4995(n4995), .n4994(n4994), 
            .n4993(n4993), .\REG.mem_5_0 (\REG.mem_5_0 ), .n4992(n4992), 
            .n4991(n4991), .n4990(n4990), .n4989(n4989), .n4988(n4988), 
            .n4987(n4987), .\REG.mem_4_10 (\REG.mem_4_10 ), .n4986(n4986), 
            .n4985(n4985), .n4984(n4984), .\REG.mem_4_7 (\REG.mem_4_7 ), 
            .n4983(n4983), .n4982(n4982), .\REG.mem_4_5 (\REG.mem_4_5 ), 
            .n4981(n4981), .n4980(n4980), .n4979(n4979), .n4978(n4978), 
            .n4977(n4977), .\REG.mem_4_0 (\REG.mem_4_0 ), .n4976(n4976), 
            .n4975(n4975), .n4974(n4974), .n4973(n4973), .n4972(n4972), 
            .n4971(n4971), .\REG.mem_3_10 (\REG.mem_3_10 ), .n4970(n4970), 
            .n4969(n4969), .\REG.mem_3_8 (\REG.mem_3_8 ), .FT_OE_N_420(FT_OE_N_420), 
            .n49(n49), .n17(n17), .n42(n42), .n10(n10), .n4968(n4968), 
            .\REG.mem_3_7 (\REG.mem_3_7 ), .n4967(n4967), .n4966(n4966), 
            .\REG.mem_3_5 (\REG.mem_3_5 ), .n4965(n4965), .n34(n34), .n4964(n4964), 
            .n4963(n4963), .n2(n2), .n4962(n4962), .n4961(n4961), .\REG.mem_3_0 (\REG.mem_3_0 ), 
            .n59(n59), .n27(n27), .n60(n60), .n28(n28), .n61(n61), 
            .n29(n29)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_dc_32_lut_gen.v(53[33] 72[34])
    
endmodule
//
// Verilog Description of module fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1
//

module fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1 (rd_addr_r, 
            \REG.mem_14_5 , \REG.mem_15_5 , \dc32_fifo_data_in[6] , dc32_fifo_almost_full, 
            FIFO_CLK_c, reset_per_frame, \REG.mem_13_5 , \REG.mem_12_5 , 
            \dc32_fifo_data_in[5] , \dc32_fifo_data_in[4] , \REG.mem_31_0 , 
            GND_net, \dc32_fifo_data_in[3] , \REG.mem_55_13 , \dc32_fifo_data_in[2] , 
            \REG.mem_38_7 , \REG.mem_39_7 , \REG.mem_36_7 , \REG.mem_37_7 , 
            \REG.mem_16_8 , \REG.mem_18_8 , \REG.mem_3_13 , \REG.mem_57_6 , 
            \dc32_fifo_data_in[1] , \REG.mem_63_11 , \dc32_fifo_data_in[0] , 
            \REG.mem_35_0 , t_rd_fifo_en_w, \REG.out_raw[0] , SLM_CLK_c, 
            \REG.mem_55_10 , n62, n30, \REG.mem_31_3 , \REG.mem_48_7 , 
            \REG.mem_50_7 , \REG.mem_55_7 , \REG.mem_48_10 , \REG.mem_50_10 , 
            wr_grey_sync_r, \wr_addr_nxt_c[5] , \REG.mem_23_8 , \REG.mem_25_5 , 
            \rd_grey_sync_r[0] , \REG.mem_25_15 , \REG.mem_14_12 , \REG.mem_15_12 , 
            DEBUG_3_c, \REG.mem_13_12 , \REG.mem_12_12 , \aempty_flag_impl.ae_flag_nxt_w , 
            dc32_fifo_almost_empty, \REG.mem_6_1 , \REG.mem_7_1 , \REG.mem_5_1 , 
            \REG.mem_4_1 , \REG.mem_57_9 , \REG.mem_35_3 , \REG.mem_46_1 , 
            \REG.mem_47_1 , \REG.mem_45_1 , \REG.mem_44_1 , \REG.mem_25_2 , 
            \dc32_fifo_data_in[15] , \dc32_fifo_data_in[14] , \dc32_fifo_data_in[13] , 
            \REG.mem_3_11 , \REG.mem_31_2 , \REG.mem_50_12 , \dc32_fifo_data_in[12] , 
            \REG.mem_6_11 , \REG.mem_7_11 , \REG.mem_5_11 , \REG.mem_4_11 , 
            \dc32_fifo_data_in[11] , \REG.mem_48_12 , \REG.mem_3_4 , \REG.mem_14_8 , 
            \REG.mem_15_8 , \REG.mem_8_14 , \REG.mem_9_14 , \dc32_fifo_data_in[10] , 
            \REG.mem_10_14 , \REG.mem_11_14 , \REG.mem_63_6 , \REG.mem_13_8 , 
            \REG.mem_12_8 , \REG.mem_14_14 , \REG.mem_15_14 , \dc32_fifo_data_in[9] , 
            \dc32_fifo_data_in[8] , \REG.mem_3_1 , \dc32_fifo_data_in[7] , 
            \REG.mem_12_14 , \REG.mem_13_14 , \REG.mem_42_8 , \REG.mem_43_8 , 
            \REG.mem_41_8 , \REG.mem_40_8 , \REG.mem_18_12 , \REG.mem_16_12 , 
            \REG.mem_31_15 , \REG.mem_38_3 , \REG.mem_39_3 , \REG.mem_37_3 , 
            \REG.mem_36_3 , \REG.mem_42_3 , \REG.mem_43_3 , \REG.mem_14_7 , 
            \REG.mem_15_7 , \REG.mem_13_7 , \REG.mem_12_7 , \REG.mem_41_3 , 
            \REG.mem_40_3 , \REG.mem_57_0 , \REG.mem_10_11 , \REG.mem_11_11 , 
            \REG.mem_9_11 , \REG.mem_8_11 , \REG.mem_63_12 , \REG.mem_55_12 , 
            \REG.mem_35_15 , \REG.mem_3_15 , \wr_addr_nxt_c[3] , \REG.mem_50_9 , 
            \REG.mem_48_9 , \REG.mem_46_8 , \REG.mem_47_8 , \REG.mem_46_3 , 
            \REG.mem_47_3 , \REG.mem_45_8 , \REG.mem_44_8 , \REG.mem_16_2 , 
            \REG.mem_10_9 , \REG.mem_11_9 , \REG.mem_45_3 , \REG.mem_44_3 , 
            \REG.mem_25_7 , \REG.mem_23_12 , \REG.mem_18_2 , \REG.mem_38_0 , 
            \REG.mem_39_0 , \REG.mem_31_13 , \REG.mem_37_0 , \REG.mem_36_0 , 
            \REG.mem_18_6 , \REG.mem_16_6 , \REG.mem_9_9 , \REG.mem_8_9 , 
            \REG.mem_50_3 , \REG.mem_48_3 , \REG.mem_42_0 , \REG.mem_43_0 , 
            \REG.mem_41_0 , \REG.mem_40_0 , \REG.mem_14_11 , \REG.mem_15_11 , 
            \REG.mem_13_11 , \REG.mem_12_11 , \REG.mem_38_5 , \REG.mem_39_5 , 
            \REG.mem_37_5 , \REG.mem_36_5 , \REG.mem_57_13 , n6121, 
            VCC_net, \fifo_data_out[2] , n6118, \fifo_data_out[1] , 
            \REG.mem_50_1 , \REG.mem_6_9 , \REG.mem_7_9 , \REG.mem_48_1 , 
            n10556, \fifo_data_out[3] , n10562, \fifo_data_out[4] , 
            \REG.mem_18_11 , \REG.mem_16_11 , \REG.mem_5_9 , \REG.mem_4_9 , 
            n10564, \fifo_data_out[5] , n10566, \fifo_data_out[6] , 
            n10568, \fifo_data_out[7] , n10570, \fifo_data_out[8] , 
            n10572, \fifo_data_out[9] , n10574, \fifo_data_out[10] , 
            n10576, \fifo_data_out[11] , \REG.mem_31_5 , n6085, \fifo_data_out[0] , 
            \REG.mem_25_12 , \REG.mem_38_13 , \REG.mem_39_13 , n10578, 
            \fifo_data_out[12] , n10580, \fifo_data_out[13] , \rd_addr_r[6] , 
            \REG.mem_6_15 , \REG.mem_7_15 , n6045, n6043, \REG.mem_5_15 , 
            \REG.mem_4_15 , \REG.mem_35_13 , n6024, n6021, \REG.mem_63_15 , 
            n6020, \REG.mem_63_14 , n6019, \REG.mem_63_13 , n6018, 
            n6017, n6016, \REG.mem_63_10 , n6015, \REG.mem_63_9 , 
            n6014, \REG.mem_63_8 , n6013, \REG.mem_63_7 , n6012, n6011, 
            \REG.mem_63_5 , n6010, \REG.mem_63_4 , n6009, \REG.mem_63_3 , 
            n6008, \REG.mem_63_2 , n6007, \REG.mem_63_1 , n6006, \REG.mem_63_0 , 
            \REG.mem_25_6 , \REG.mem_37_13 , \REG.mem_36_13 , \REG.mem_57_4 , 
            \REG.mem_18_7 , \REG.mem_16_7 , \REG.mem_38_15 , \REG.mem_39_15 , 
            \REG.mem_23_11 , \REG.mem_37_15 , \REG.mem_36_15 , \REG.mem_25_11 , 
            \REG.mem_57_12 , \REG.mem_40_14 , \REG.mem_41_14 , n5953, 
            rp_sync1_r, \REG.mem_42_14 , \REG.mem_43_14 , \REG.mem_46_14 , 
            \REG.mem_47_14 , n5952, n5951, n5950, n5949, n5948, 
            n5947, n5946, n5945, \REG.mem_55_9 , \REG.mem_44_14 , 
            \REG.mem_45_14 , \REG.mem_10_7 , \REG.mem_11_7 , n5928, 
            n5927, n5926, n5924, n5923, n5921, \REG.mem_9_7 , \REG.mem_8_7 , 
            \REG.mem_40_4 , \REG.mem_41_4 , \REG.mem_42_4 , \REG.mem_43_4 , 
            \REG.mem_46_4 , \REG.mem_47_4 , \REG.mem_44_4 , \REG.mem_45_4 , 
            n5901, \REG.mem_57_15 , n5900, \REG.mem_57_14 , n5899, 
            n5898, n5897, \REG.mem_57_11 , n5896, \REG.mem_57_10 , 
            n5895, n5894, \REG.mem_57_8 , n5893, \REG.mem_57_7 , n5892, 
            n5891, \REG.mem_57_5 , n5890, n5889, \REG.mem_57_3 , n5888, 
            \REG.mem_57_2 , n5887, \REG.mem_57_1 , \REG.mem_18_1 , \REG.mem_16_1 , 
            n5885, \REG.mem_35_8 , \REG.mem_38_8 , \REG.mem_39_8 , \REG.mem_36_8 , 
            \REG.mem_37_8 , n5864, wp_sync1_r, n5863, n5862, n5861, 
            n5860, n5859, n5858, \REG.mem_55_15 , n5857, \REG.mem_55_14 , 
            n5856, n5855, n5854, \REG.mem_55_11 , n5853, \rd_sig_diff0_w[0] , 
            n5852, n5851, \REG.mem_55_8 , n5850, n5849, \REG.mem_55_6 , 
            n5848, \REG.mem_55_5 , n5847, \REG.mem_55_4 , n5846, \REG.mem_55_3 , 
            n5845, \REG.mem_55_2 , n5844, \REG.mem_55_1 , n5843, \REG.mem_55_0 , 
            n5842, n5841, n5839, n5838, n5837, \REG.mem_16_15 , 
            \REG.mem_18_15 , \REG.mem_23_15 , n5836, \REG.mem_25_4 , 
            \REG.mem_35_2 , \REG.mem_31_4 , \REG.mem_38_2 , \REG.mem_39_2 , 
            \REG.mem_36_2 , \REG.mem_37_2 , \REG.mem_10_15 , \REG.mem_11_15 , 
            \REG.mem_48_2 , \REG.mem_50_2 , \REG.mem_8_4 , \REG.mem_9_4 , 
            \REG.mem_10_4 , \REG.mem_11_4 , n5771, \REG.mem_50_15 , 
            n5770, \REG.mem_50_14 , n5769, \REG.mem_50_13 , n5768, 
            n5767, \REG.mem_50_11 , n5766, n5765, n5764, \REG.mem_50_8 , 
            n5763, n5762, \REG.mem_50_6 , n5761, \REG.mem_50_5 , n5760, 
            \REG.mem_50_4 , n5759, n5758, n5757, \REG.mem_14_4 , \REG.mem_15_4 , 
            n10873, \REG.mem_12_4 , \REG.mem_13_4 , n10582, \fifo_data_out[14] , 
            n10588, \fifo_data_out[15] , n5753, \REG.mem_50_0 , \REG.mem_3_14 , 
            \REG.mem_6_14 , \REG.mem_7_14 , \REG.mem_4_14 , \REG.mem_5_14 , 
            n5736, \REG.mem_48_15 , n5735, \REG.mem_48_14 , n5734, 
            \REG.mem_48_13 , n5733, n5732, \REG.mem_48_11 , n5731, 
            n5730, n5729, \REG.mem_48_8 , n5728, n5727, \REG.mem_48_6 , 
            n5726, \REG.mem_48_5 , n5725, \REG.mem_48_4 , n5724, n10877, 
            \REG.mem_9_15 , \REG.mem_8_15 , \REG.mem_31_7 , n5723, n5722, 
            n5721, \REG.mem_48_0 , n5720, \REG.mem_47_15 , n5719, 
            n5718, \REG.mem_47_13 , n5717, \REG.mem_47_12 , n5716, 
            \REG.mem_47_11 , n5715, \REG.mem_47_10 , n5714, \REG.mem_47_9 , 
            n5713, n5712, \REG.mem_47_7 , n5711, \REG.mem_47_6 , n5710, 
            \REG.mem_47_5 , n5709, n5708, n5707, \REG.mem_47_2 , n5706, 
            n5705, \REG.mem_47_0 , n5704, \REG.mem_46_15 , n5703, 
            \REG.mem_31_12 , n5702, \REG.mem_46_13 , n5701, \REG.mem_46_12 , 
            n5700, \REG.mem_46_11 , n5699, \REG.mem_46_10 , n5698, 
            \REG.mem_46_9 , n5697, n5696, \REG.mem_46_7 , n5695, \REG.mem_46_6 , 
            n5694, \REG.mem_46_5 , n5693, n5692, n5691, \REG.mem_46_2 , 
            n5690, n5689, \REG.mem_46_0 , n5688, \REG.mem_45_15 , 
            n5687, n5686, \REG.mem_45_13 , n5685, \REG.mem_45_12 , 
            n5684, \REG.mem_45_11 , n5683, \REG.mem_45_10 , n5682, 
            \REG.mem_45_9 , n5681, n5680, \REG.mem_45_7 , n5679, \REG.mem_45_6 , 
            n5678, \REG.mem_45_5 , \REG.mem_38_6 , \REG.mem_39_6 , \REG.mem_37_6 , 
            \REG.mem_36_6 , n5677, \REG.mem_31_11 , n5676, \REG.mem_42_5 , 
            \REG.mem_43_5 , n5675, \REG.mem_45_2 , n5674, n5673, \REG.mem_45_0 , 
            n5671, \REG.mem_44_15 , n5670, n5669, \REG.mem_44_13 , 
            n5668, \REG.mem_44_12 , n5666, \REG.mem_44_11 , n5665, 
            \REG.mem_44_10 , n5664, \REG.mem_44_9 , n5662, n5661, 
            \REG.mem_44_7 , n5660, \REG.mem_44_6 , n5659, \REG.mem_44_5 , 
            n5658, n5657, n5656, \REG.mem_44_2 , n5655, n5654, \REG.mem_44_0 , 
            n5653, \REG.mem_43_15 , n5652, n5651, \REG.mem_43_13 , 
            n5650, \REG.mem_43_12 , n5649, \REG.mem_43_11 , n5648, 
            \REG.mem_43_10 , n5647, \REG.mem_43_9 , n5646, n5645, 
            \REG.mem_43_7 , n5644, \REG.mem_43_6 , \REG.mem_41_5 , \REG.mem_40_5 , 
            \REG.mem_23_1 , \rd_addr_p1_w[0] , \REG.mem_35_11 , n5643, 
            n5642, n5641, n5640, \REG.mem_43_2 , n5639, \REG.mem_43_1 , 
            n5638, n5637, \REG.mem_42_15 , n5636, n5635, \REG.mem_42_13 , 
            n5634, \REG.mem_42_12 , n5633, \REG.mem_42_11 , n5632, 
            \REG.mem_42_10 , n5631, \REG.mem_42_9 , n5630, n5629, 
            \REG.mem_42_7 , n4916, \REG.mem_31_6 , \REG.mem_23_2 , \REG.mem_38_11 , 
            \REG.mem_39_11 , \REG.mem_37_11 , \REG.mem_36_11 , n5628, 
            \REG.mem_42_6 , n5627, n5626, n5625, n5624, \REG.mem_42_2 , 
            n5623, \REG.mem_42_1 , n5622, n5621, \REG.mem_41_15 , 
            n5620, n5619, \REG.mem_41_13 , n5618, \REG.mem_41_12 , 
            n5617, \REG.mem_41_11 , n5616, \REG.mem_41_10 , n5615, 
            \REG.mem_41_9 , n5614, n5613, \REG.mem_41_7 , \REG.mem_3_2 , 
            n5612, \REG.mem_41_6 , n5611, n5610, n5609, n5608, \REG.mem_41_2 , 
            n5607, \REG.mem_41_1 , n5606, n5605, \REG.mem_40_15 , 
            n5604, n5603, \REG.mem_40_13 , n5602, \REG.mem_40_12 , 
            n5601, \REG.mem_40_11 , n5600, \REG.mem_40_10 , n5599, 
            \REG.mem_40_9 , n5598, n5597, \REG.mem_40_7 , \REG.mem_25_9 , 
            n4904, n4903, n4901, n4899, n5596, \REG.mem_40_6 , n5595, 
            n5594, n5593, n5592, \REG.mem_40_2 , n5591, \REG.mem_40_1 , 
            n5590, n5589, n5588, \REG.mem_39_14 , n5587, n5586, 
            \REG.mem_39_12 , n5585, n5584, \REG.mem_39_10 , n5583, 
            \REG.mem_39_9 , n5582, n5581, n4898, \REG.mem_14_1 , \REG.mem_15_1 , 
            DEBUG_5_c, \REG.mem_13_1 , \REG.mem_12_1 , \REG.mem_3_3 , 
            n5580, n5579, n5578, \REG.mem_39_4 , n5577, n5576, n5575, 
            \REG.mem_39_1 , n5573, n5572, n5571, \REG.mem_38_14 , 
            n5570, n5569, \REG.mem_38_12 , n5568, n5567, \REG.mem_38_10 , 
            n5566, \REG.mem_38_9 , n5565, n5564, n5563, n5562, n5561, 
            \REG.mem_38_4 , n5560, n5559, n5558, \REG.mem_38_1 , n5556, 
            n5555, n5554, \REG.mem_37_14 , n5553, n5552, \REG.mem_37_12 , 
            n5551, n5550, \REG.mem_37_10 , n5549, \REG.mem_37_9 , 
            \REG.mem_25_13 , \REG.out_raw[15] , \REG.out_raw[14] , \REG.out_raw[13] , 
            \REG.out_raw[12] , \REG.out_raw[11] , n5548, n5547, n5546, 
            n5545, n5544, \REG.mem_37_4 , n5543, n5542, n5541, \REG.mem_37_1 , 
            n5540, \REG.out_raw[10] , \REG.out_raw[9] , \REG.out_raw[8] , 
            \REG.out_raw[7] , \REG.out_raw[6] , \REG.out_raw[5] , \REG.out_raw[4] , 
            \REG.out_raw[3] , \REG.out_raw[2] , \REG.out_raw[1] , n5526, 
            n5525, \REG.mem_36_14 , n5524, n5523, \REG.mem_36_12 , 
            n5522, n5521, \REG.mem_36_10 , n5520, \REG.mem_36_9 , 
            n5519, n5518, n5517, n5516, \rd_sig_diff0_w[2] , n5515, 
            \REG.mem_36_4 , n5514, n5513, n5512, \REG.mem_36_1 , n5511, 
            n5507, n5506, \REG.mem_35_14 , n5505, n5504, \REG.mem_35_12 , 
            n5503, n5502, \REG.mem_35_10 , n5501, \REG.mem_35_9 , 
            n5500, \rd_sig_diff0_w[1] , n5499, \REG.mem_35_7 , n5498, 
            \REG.mem_35_6 , n5497, \REG.mem_35_5 , n5496, \REG.mem_35_4 , 
            n5495, n5494, n5493, \REG.mem_35_1 , n5492, \REG.mem_6_3 , 
            \REG.mem_7_3 , \REG.mem_5_3 , \REG.mem_4_3 , n5441, n5440, 
            \REG.mem_31_14 , n5439, n5438, n5437, \REG.mem_25_1 , 
            n5436, \REG.mem_31_10 , n58, n5435, \REG.mem_31_9 , n5434, 
            \REG.mem_31_8 , n5433, n5432, n5431, n5430, n5429, n5428, 
            n5427, \REG.mem_31_1 , n5426, n26, DEBUG_1_c_c, write_to_dc32_fifo_latched_N_425, 
            n5345, n5344, \REG.mem_25_14 , n5343, n5342, n5341, 
            n5340, \REG.mem_25_10 , n5339, n5338, \REG.mem_25_8 , 
            n5337, n5336, n5335, n5334, n5333, \REG.mem_25_3 , n5332, 
            n5331, n5330, \REG.mem_25_0 , \REG.mem_14_15 , \REG.mem_15_15 , 
            \REG.mem_6_13 , \REG.mem_7_13 , n5306, n5305, \REG.mem_23_14 , 
            n5304, \REG.mem_23_13 , n5303, n5302, n5301, \REG.mem_23_10 , 
            n5300, \REG.mem_23_9 , n5299, n5298, \REG.mem_23_7 , n5297, 
            \REG.mem_23_6 , n5296, \REG.mem_23_5 , n5295, \REG.mem_23_4 , 
            n5294, \REG.mem_23_3 , n5293, n5292, n5290, \REG.mem_23_0 , 
            \rd_grey_sync_r[5] , \REG.mem_5_13 , \REG.mem_4_13 , \rd_grey_sync_r[4] , 
            \rd_grey_sync_r[3] , \rd_grey_sync_r[2] , \rd_grey_sync_r[1] , 
            \REG.mem_13_15 , \REG.mem_12_15 , n51, n19, \wr_addr_nxt_c[1] , 
            \REG.mem_10_0 , \REG.mem_11_0 , \REG.mem_10_3 , \REG.mem_11_3 , 
            n5224, n5223, \REG.mem_18_14 , n5222, \REG.mem_18_13 , 
            n5221, n5220, \REG.mem_9_3 , \REG.mem_8_3 , \REG.mem_9_0 , 
            \REG.mem_8_0 , \REG.mem_10_13 , \REG.mem_11_13 , n52, \REG.mem_9_13 , 
            \REG.mem_8_13 , n20, n5219, \REG.mem_18_10 , n5218, \REG.mem_18_9 , 
            n5217, n5216, n5215, n5214, \REG.mem_18_5 , n5213, \REG.mem_18_4 , 
            n5212, \REG.mem_18_3 , n5211, n5210, n5209, \REG.mem_18_0 , 
            \REG.mem_14_13 , \REG.mem_15_13 , \REG.mem_13_13 , \REG.mem_12_13 , 
            \REG.mem_6_4 , \REG.mem_7_4 , \REG.mem_5_4 , \REG.mem_4_4 , 
            get_next_word, n5188, n5186, \REG.mem_16_14 , n5185, \REG.mem_16_13 , 
            \REG.mem_6_8 , \REG.mem_7_8 , \REG.mem_3_6 , n5184, \REG.mem_5_8 , 
            \REG.mem_4_8 , \REG.mem_6_2 , \REG.mem_7_2 , \REG.mem_5_2 , 
            \REG.mem_4_2 , rd_fifo_en_w, n5183, n5182, \REG.mem_16_10 , 
            n5181, \REG.mem_16_9 , n5180, n5179, n5178, n5177, \REG.mem_16_5 , 
            n5176, \REG.mem_16_4 , \REG.mem_3_12 , n5175, \REG.mem_16_3 , 
            n5174, n5173, n5172, \REG.mem_16_0 , n5169, n5168, n5167, 
            n47, n5166, n15, n5165, n5164, \REG.mem_15_10 , n5163, 
            \REG.mem_15_9 , n5162, n5161, n5160, \REG.mem_15_6 , n5159, 
            n5158, n5157, \REG.mem_15_3 , n5156, \REG.mem_15_2 , n5155, 
            n5154, \REG.mem_15_0 , n5153, n5152, \REG.mem_6_6 , \REG.mem_7_6 , 
            n5151, n5150, n5149, n5148, \REG.mem_14_10 , n5147, 
            \REG.mem_14_9 , n5146, n5145, n5144, \REG.mem_14_6 , \REG.mem_4_6 , 
            \REG.mem_5_6 , n5143, n5142, n5141, \REG.mem_14_3 , n5140, 
            \REG.mem_14_2 , n5139, n5138, \REG.mem_14_0 , n5137, n5136, 
            n5135, n5134, n5133, n5132, \REG.mem_13_10 , \REG.mem_13_9 , 
            \REG.mem_12_9 , n5131, n5130, n5129, n5128, \REG.mem_13_6 , 
            n5127, n5126, n5125, \REG.mem_13_3 , n5124, \REG.mem_13_2 , 
            n5123, \REG.mem_10_8 , \REG.mem_11_8 , n5122, \REG.mem_13_0 , 
            n5121, n5120, n5119, n5118, \REG.mem_3_9 , \REG.mem_9_8 , 
            \REG.mem_8_8 , n5117, \REG.mem_8_6 , \REG.mem_9_6 , n5116, 
            \REG.mem_12_10 , \REG.mem_10_6 , \REG.mem_11_6 , n53, n21, 
            n5115, n5114, n5113, n5112, \REG.mem_12_6 , n50, n5111, 
            n18, \REG.mem_6_12 , \REG.mem_7_12 , n5110, n5109, \REG.mem_12_3 , 
            n5108, \REG.mem_12_2 , \REG.mem_4_12 , \REG.mem_5_12 , \REG.mem_10_2 , 
            \REG.mem_11_2 , n5107, \REG.mem_9_2 , \REG.mem_8_2 , n54, 
            n22, n5106, \REG.mem_12_0 , \rd_addr_nxt_c_6__N_498[3] , 
            n5105, n5104, n5103, n5102, \REG.mem_11_12 , n5101, 
            n5100, \REG.mem_11_10 , n5099, n5098, n5097, n5096, 
            n5095, \REG.mem_11_5 , n5094, n5093, n5092, n5091, \REG.mem_11_1 , 
            n5090, n5089, n5088, \rd_addr_nxt_c_6__N_498[5] , n5087, 
            n5086, \REG.mem_10_12 , n5085, n5084, \REG.mem_10_10 , 
            n5083, n5082, n5081, n5080, n5079, \REG.mem_10_5 , \REG.mem_10_1 , 
            \REG.mem_9_1 , \REG.mem_8_1 , \rd_addr_nxt_c_6__N_498[2] , 
            n56, n24, n5078, n55, n23, n5077, n40, n8, n5076, 
            n5075, n5074, n5073, n5072, n5071, n5070, \REG.mem_9_12 , 
            n5069, n5068, \REG.mem_9_10 , n5067, n5066, n5065, n57, 
            n5064, n25, n5063, \REG.mem_9_5 , n5062, n5061, n5060, 
            n5059, n5057, n5056, n5055, n5054, n5053, \REG.mem_8_12 , 
            n5052, n5051, \REG.mem_8_10 , n5050, n5049, n5048, n5047, 
            n5046, \REG.mem_8_5 , n5045, n5044, n5043, n5042, n5041, 
            n5040, n5039, n5038, n5037, n5036, n5035, \REG.mem_7_10 , 
            n5034, n5033, n5032, \REG.mem_7_7 , n5031, n5030, \REG.mem_7_5 , 
            n5029, n5028, n5027, n5026, n5025, \REG.mem_7_0 , n5024, 
            n5023, n5022, n5021, n5020, n5019, \REG.mem_6_10 , n5018, 
            n5017, n5016, \REG.mem_6_7 , n5015, n5014, \REG.mem_6_5 , 
            n5013, n5012, n5011, n5010, n5009, \REG.mem_6_0 , n5008, 
            n5007, n5006, n5005, n5004, n5003, \REG.mem_5_10 , n5002, 
            n5001, n5000, \REG.mem_5_7 , n4999, n4998, \REG.mem_5_5 , 
            n4997, n4996, n4995, n4994, n4993, \REG.mem_5_0 , n4992, 
            n4991, n4990, n4989, n4988, n4987, \REG.mem_4_10 , n4986, 
            n4985, n4984, \REG.mem_4_7 , n4983, n4982, \REG.mem_4_5 , 
            n4981, n4980, n4979, n4978, n4977, \REG.mem_4_0 , n4976, 
            n4975, n4974, n4973, n4972, n4971, \REG.mem_3_10 , n4970, 
            n4969, \REG.mem_3_8 , FT_OE_N_420, n49, n17, n42, n10, 
            n4968, \REG.mem_3_7 , n4967, n4966, \REG.mem_3_5 , n4965, 
            n34, n4964, n4963, n2, n4962, n4961, \REG.mem_3_0 , 
            n59, n27, n60, n28, n61, n29) /* synthesis syn_module_defined=1 */ ;
    output [6:0]rd_addr_r;
    output \REG.mem_14_5 ;
    output \REG.mem_15_5 ;
    input \dc32_fifo_data_in[6] ;
    output dc32_fifo_almost_full;
    input FIFO_CLK_c;
    input reset_per_frame;
    output \REG.mem_13_5 ;
    output \REG.mem_12_5 ;
    input \dc32_fifo_data_in[5] ;
    input \dc32_fifo_data_in[4] ;
    output \REG.mem_31_0 ;
    input GND_net;
    input \dc32_fifo_data_in[3] ;
    output \REG.mem_55_13 ;
    input \dc32_fifo_data_in[2] ;
    output \REG.mem_38_7 ;
    output \REG.mem_39_7 ;
    output \REG.mem_36_7 ;
    output \REG.mem_37_7 ;
    output \REG.mem_16_8 ;
    output \REG.mem_18_8 ;
    output \REG.mem_3_13 ;
    output \REG.mem_57_6 ;
    input \dc32_fifo_data_in[1] ;
    output \REG.mem_63_11 ;
    input \dc32_fifo_data_in[0] ;
    output \REG.mem_35_0 ;
    output t_rd_fifo_en_w;
    output \REG.out_raw[0] ;
    input SLM_CLK_c;
    output \REG.mem_55_10 ;
    output n62;
    output n30;
    output \REG.mem_31_3 ;
    output \REG.mem_48_7 ;
    output \REG.mem_50_7 ;
    output \REG.mem_55_7 ;
    output \REG.mem_48_10 ;
    output \REG.mem_50_10 ;
    output [6:0]wr_grey_sync_r;
    output \wr_addr_nxt_c[5] ;
    output \REG.mem_23_8 ;
    output \REG.mem_25_5 ;
    output \rd_grey_sync_r[0] ;
    output \REG.mem_25_15 ;
    output \REG.mem_14_12 ;
    output \REG.mem_15_12 ;
    output DEBUG_3_c;
    output \REG.mem_13_12 ;
    output \REG.mem_12_12 ;
    input \aempty_flag_impl.ae_flag_nxt_w ;
    output dc32_fifo_almost_empty;
    output \REG.mem_6_1 ;
    output \REG.mem_7_1 ;
    output \REG.mem_5_1 ;
    output \REG.mem_4_1 ;
    output \REG.mem_57_9 ;
    output \REG.mem_35_3 ;
    output \REG.mem_46_1 ;
    output \REG.mem_47_1 ;
    output \REG.mem_45_1 ;
    output \REG.mem_44_1 ;
    output \REG.mem_25_2 ;
    input \dc32_fifo_data_in[15] ;
    input \dc32_fifo_data_in[14] ;
    input \dc32_fifo_data_in[13] ;
    output \REG.mem_3_11 ;
    output \REG.mem_31_2 ;
    output \REG.mem_50_12 ;
    input \dc32_fifo_data_in[12] ;
    output \REG.mem_6_11 ;
    output \REG.mem_7_11 ;
    output \REG.mem_5_11 ;
    output \REG.mem_4_11 ;
    input \dc32_fifo_data_in[11] ;
    output \REG.mem_48_12 ;
    output \REG.mem_3_4 ;
    output \REG.mem_14_8 ;
    output \REG.mem_15_8 ;
    output \REG.mem_8_14 ;
    output \REG.mem_9_14 ;
    input \dc32_fifo_data_in[10] ;
    output \REG.mem_10_14 ;
    output \REG.mem_11_14 ;
    output \REG.mem_63_6 ;
    output \REG.mem_13_8 ;
    output \REG.mem_12_8 ;
    output \REG.mem_14_14 ;
    output \REG.mem_15_14 ;
    input \dc32_fifo_data_in[9] ;
    input \dc32_fifo_data_in[8] ;
    output \REG.mem_3_1 ;
    input \dc32_fifo_data_in[7] ;
    output \REG.mem_12_14 ;
    output \REG.mem_13_14 ;
    output \REG.mem_42_8 ;
    output \REG.mem_43_8 ;
    output \REG.mem_41_8 ;
    output \REG.mem_40_8 ;
    output \REG.mem_18_12 ;
    output \REG.mem_16_12 ;
    output \REG.mem_31_15 ;
    output \REG.mem_38_3 ;
    output \REG.mem_39_3 ;
    output \REG.mem_37_3 ;
    output \REG.mem_36_3 ;
    output \REG.mem_42_3 ;
    output \REG.mem_43_3 ;
    output \REG.mem_14_7 ;
    output \REG.mem_15_7 ;
    output \REG.mem_13_7 ;
    output \REG.mem_12_7 ;
    output \REG.mem_41_3 ;
    output \REG.mem_40_3 ;
    output \REG.mem_57_0 ;
    output \REG.mem_10_11 ;
    output \REG.mem_11_11 ;
    output \REG.mem_9_11 ;
    output \REG.mem_8_11 ;
    output \REG.mem_63_12 ;
    output \REG.mem_55_12 ;
    output \REG.mem_35_15 ;
    output \REG.mem_3_15 ;
    output \wr_addr_nxt_c[3] ;
    output \REG.mem_50_9 ;
    output \REG.mem_48_9 ;
    output \REG.mem_46_8 ;
    output \REG.mem_47_8 ;
    output \REG.mem_46_3 ;
    output \REG.mem_47_3 ;
    output \REG.mem_45_8 ;
    output \REG.mem_44_8 ;
    output \REG.mem_16_2 ;
    output \REG.mem_10_9 ;
    output \REG.mem_11_9 ;
    output \REG.mem_45_3 ;
    output \REG.mem_44_3 ;
    output \REG.mem_25_7 ;
    output \REG.mem_23_12 ;
    output \REG.mem_18_2 ;
    output \REG.mem_38_0 ;
    output \REG.mem_39_0 ;
    output \REG.mem_31_13 ;
    output \REG.mem_37_0 ;
    output \REG.mem_36_0 ;
    output \REG.mem_18_6 ;
    output \REG.mem_16_6 ;
    output \REG.mem_9_9 ;
    output \REG.mem_8_9 ;
    output \REG.mem_50_3 ;
    output \REG.mem_48_3 ;
    output \REG.mem_42_0 ;
    output \REG.mem_43_0 ;
    output \REG.mem_41_0 ;
    output \REG.mem_40_0 ;
    output \REG.mem_14_11 ;
    output \REG.mem_15_11 ;
    output \REG.mem_13_11 ;
    output \REG.mem_12_11 ;
    output \REG.mem_38_5 ;
    output \REG.mem_39_5 ;
    output \REG.mem_37_5 ;
    output \REG.mem_36_5 ;
    output \REG.mem_57_13 ;
    input n6121;
    input VCC_net;
    output \fifo_data_out[2] ;
    input n6118;
    output \fifo_data_out[1] ;
    output \REG.mem_50_1 ;
    output \REG.mem_6_9 ;
    output \REG.mem_7_9 ;
    output \REG.mem_48_1 ;
    input n10556;
    output \fifo_data_out[3] ;
    input n10562;
    output \fifo_data_out[4] ;
    output \REG.mem_18_11 ;
    output \REG.mem_16_11 ;
    output \REG.mem_5_9 ;
    output \REG.mem_4_9 ;
    input n10564;
    output \fifo_data_out[5] ;
    input n10566;
    output \fifo_data_out[6] ;
    input n10568;
    output \fifo_data_out[7] ;
    input n10570;
    output \fifo_data_out[8] ;
    input n10572;
    output \fifo_data_out[9] ;
    input n10574;
    output \fifo_data_out[10] ;
    input n10576;
    output \fifo_data_out[11] ;
    output \REG.mem_31_5 ;
    input n6085;
    output \fifo_data_out[0] ;
    output \REG.mem_25_12 ;
    output \REG.mem_38_13 ;
    output \REG.mem_39_13 ;
    input n10578;
    output \fifo_data_out[12] ;
    input n10580;
    output \fifo_data_out[13] ;
    output \rd_addr_r[6] ;
    output \REG.mem_6_15 ;
    output \REG.mem_7_15 ;
    input n6045;
    input n6043;
    output \REG.mem_5_15 ;
    output \REG.mem_4_15 ;
    output \REG.mem_35_13 ;
    input n6024;
    input n6021;
    output \REG.mem_63_15 ;
    input n6020;
    output \REG.mem_63_14 ;
    input n6019;
    output \REG.mem_63_13 ;
    input n6018;
    input n6017;
    input n6016;
    output \REG.mem_63_10 ;
    input n6015;
    output \REG.mem_63_9 ;
    input n6014;
    output \REG.mem_63_8 ;
    input n6013;
    output \REG.mem_63_7 ;
    input n6012;
    input n6011;
    output \REG.mem_63_5 ;
    input n6010;
    output \REG.mem_63_4 ;
    input n6009;
    output \REG.mem_63_3 ;
    input n6008;
    output \REG.mem_63_2 ;
    input n6007;
    output \REG.mem_63_1 ;
    input n6006;
    output \REG.mem_63_0 ;
    output \REG.mem_25_6 ;
    output \REG.mem_37_13 ;
    output \REG.mem_36_13 ;
    output \REG.mem_57_4 ;
    output \REG.mem_18_7 ;
    output \REG.mem_16_7 ;
    output \REG.mem_38_15 ;
    output \REG.mem_39_15 ;
    output \REG.mem_23_11 ;
    output \REG.mem_37_15 ;
    output \REG.mem_36_15 ;
    output \REG.mem_25_11 ;
    output \REG.mem_57_12 ;
    output \REG.mem_40_14 ;
    output \REG.mem_41_14 ;
    input n5953;
    output [6:0]rp_sync1_r;
    output \REG.mem_42_14 ;
    output \REG.mem_43_14 ;
    output \REG.mem_46_14 ;
    output \REG.mem_47_14 ;
    input n5952;
    input n5951;
    input n5950;
    input n5949;
    input n5948;
    input n5947;
    input n5946;
    input n5945;
    output \REG.mem_55_9 ;
    output \REG.mem_44_14 ;
    output \REG.mem_45_14 ;
    output \REG.mem_10_7 ;
    output \REG.mem_11_7 ;
    input n5928;
    input n5927;
    input n5926;
    input n5924;
    input n5923;
    input n5921;
    output \REG.mem_9_7 ;
    output \REG.mem_8_7 ;
    output \REG.mem_40_4 ;
    output \REG.mem_41_4 ;
    output \REG.mem_42_4 ;
    output \REG.mem_43_4 ;
    output \REG.mem_46_4 ;
    output \REG.mem_47_4 ;
    output \REG.mem_44_4 ;
    output \REG.mem_45_4 ;
    input n5901;
    output \REG.mem_57_15 ;
    input n5900;
    output \REG.mem_57_14 ;
    input n5899;
    input n5898;
    input n5897;
    output \REG.mem_57_11 ;
    input n5896;
    output \REG.mem_57_10 ;
    input n5895;
    input n5894;
    output \REG.mem_57_8 ;
    input n5893;
    output \REG.mem_57_7 ;
    input n5892;
    input n5891;
    output \REG.mem_57_5 ;
    input n5890;
    input n5889;
    output \REG.mem_57_3 ;
    input n5888;
    output \REG.mem_57_2 ;
    input n5887;
    output \REG.mem_57_1 ;
    output \REG.mem_18_1 ;
    output \REG.mem_16_1 ;
    input n5885;
    output \REG.mem_35_8 ;
    output \REG.mem_38_8 ;
    output \REG.mem_39_8 ;
    output \REG.mem_36_8 ;
    output \REG.mem_37_8 ;
    input n5864;
    output [6:0]wp_sync1_r;
    input n5863;
    input n5862;
    input n5861;
    input n5860;
    input n5859;
    input n5858;
    output \REG.mem_55_15 ;
    input n5857;
    output \REG.mem_55_14 ;
    input n5856;
    input n5855;
    input n5854;
    output \REG.mem_55_11 ;
    input n5853;
    output \rd_sig_diff0_w[0] ;
    input n5852;
    input n5851;
    output \REG.mem_55_8 ;
    input n5850;
    input n5849;
    output \REG.mem_55_6 ;
    input n5848;
    output \REG.mem_55_5 ;
    input n5847;
    output \REG.mem_55_4 ;
    input n5846;
    output \REG.mem_55_3 ;
    input n5845;
    output \REG.mem_55_2 ;
    input n5844;
    output \REG.mem_55_1 ;
    input n5843;
    output \REG.mem_55_0 ;
    input n5842;
    input n5841;
    input n5839;
    input n5838;
    input n5837;
    output \REG.mem_16_15 ;
    output \REG.mem_18_15 ;
    output \REG.mem_23_15 ;
    input n5836;
    output \REG.mem_25_4 ;
    output \REG.mem_35_2 ;
    output \REG.mem_31_4 ;
    output \REG.mem_38_2 ;
    output \REG.mem_39_2 ;
    output \REG.mem_36_2 ;
    output \REG.mem_37_2 ;
    output \REG.mem_10_15 ;
    output \REG.mem_11_15 ;
    output \REG.mem_48_2 ;
    output \REG.mem_50_2 ;
    output \REG.mem_8_4 ;
    output \REG.mem_9_4 ;
    output \REG.mem_10_4 ;
    output \REG.mem_11_4 ;
    input n5771;
    output \REG.mem_50_15 ;
    input n5770;
    output \REG.mem_50_14 ;
    input n5769;
    output \REG.mem_50_13 ;
    input n5768;
    input n5767;
    output \REG.mem_50_11 ;
    input n5766;
    input n5765;
    input n5764;
    output \REG.mem_50_8 ;
    input n5763;
    input n5762;
    output \REG.mem_50_6 ;
    input n5761;
    output \REG.mem_50_5 ;
    input n5760;
    output \REG.mem_50_4 ;
    input n5759;
    input n5758;
    input n5757;
    output \REG.mem_14_4 ;
    output \REG.mem_15_4 ;
    output n10873;
    output \REG.mem_12_4 ;
    output \REG.mem_13_4 ;
    input n10582;
    output \fifo_data_out[14] ;
    input n10588;
    output \fifo_data_out[15] ;
    input n5753;
    output \REG.mem_50_0 ;
    output \REG.mem_3_14 ;
    output \REG.mem_6_14 ;
    output \REG.mem_7_14 ;
    output \REG.mem_4_14 ;
    output \REG.mem_5_14 ;
    input n5736;
    output \REG.mem_48_15 ;
    input n5735;
    output \REG.mem_48_14 ;
    input n5734;
    output \REG.mem_48_13 ;
    input n5733;
    input n5732;
    output \REG.mem_48_11 ;
    input n5731;
    input n5730;
    input n5729;
    output \REG.mem_48_8 ;
    input n5728;
    input n5727;
    output \REG.mem_48_6 ;
    input n5726;
    output \REG.mem_48_5 ;
    input n5725;
    output \REG.mem_48_4 ;
    input n5724;
    output n10877;
    output \REG.mem_9_15 ;
    output \REG.mem_8_15 ;
    output \REG.mem_31_7 ;
    input n5723;
    input n5722;
    input n5721;
    output \REG.mem_48_0 ;
    input n5720;
    output \REG.mem_47_15 ;
    input n5719;
    input n5718;
    output \REG.mem_47_13 ;
    input n5717;
    output \REG.mem_47_12 ;
    input n5716;
    output \REG.mem_47_11 ;
    input n5715;
    output \REG.mem_47_10 ;
    input n5714;
    output \REG.mem_47_9 ;
    input n5713;
    input n5712;
    output \REG.mem_47_7 ;
    input n5711;
    output \REG.mem_47_6 ;
    input n5710;
    output \REG.mem_47_5 ;
    input n5709;
    input n5708;
    input n5707;
    output \REG.mem_47_2 ;
    input n5706;
    input n5705;
    output \REG.mem_47_0 ;
    input n5704;
    output \REG.mem_46_15 ;
    input n5703;
    output \REG.mem_31_12 ;
    input n5702;
    output \REG.mem_46_13 ;
    input n5701;
    output \REG.mem_46_12 ;
    input n5700;
    output \REG.mem_46_11 ;
    input n5699;
    output \REG.mem_46_10 ;
    input n5698;
    output \REG.mem_46_9 ;
    input n5697;
    input n5696;
    output \REG.mem_46_7 ;
    input n5695;
    output \REG.mem_46_6 ;
    input n5694;
    output \REG.mem_46_5 ;
    input n5693;
    input n5692;
    input n5691;
    output \REG.mem_46_2 ;
    input n5690;
    input n5689;
    output \REG.mem_46_0 ;
    input n5688;
    output \REG.mem_45_15 ;
    input n5687;
    input n5686;
    output \REG.mem_45_13 ;
    input n5685;
    output \REG.mem_45_12 ;
    input n5684;
    output \REG.mem_45_11 ;
    input n5683;
    output \REG.mem_45_10 ;
    input n5682;
    output \REG.mem_45_9 ;
    input n5681;
    input n5680;
    output \REG.mem_45_7 ;
    input n5679;
    output \REG.mem_45_6 ;
    input n5678;
    output \REG.mem_45_5 ;
    output \REG.mem_38_6 ;
    output \REG.mem_39_6 ;
    output \REG.mem_37_6 ;
    output \REG.mem_36_6 ;
    input n5677;
    output \REG.mem_31_11 ;
    input n5676;
    output \REG.mem_42_5 ;
    output \REG.mem_43_5 ;
    input n5675;
    output \REG.mem_45_2 ;
    input n5674;
    input n5673;
    output \REG.mem_45_0 ;
    input n5671;
    output \REG.mem_44_15 ;
    input n5670;
    input n5669;
    output \REG.mem_44_13 ;
    input n5668;
    output \REG.mem_44_12 ;
    input n5666;
    output \REG.mem_44_11 ;
    input n5665;
    output \REG.mem_44_10 ;
    input n5664;
    output \REG.mem_44_9 ;
    input n5662;
    input n5661;
    output \REG.mem_44_7 ;
    input n5660;
    output \REG.mem_44_6 ;
    input n5659;
    output \REG.mem_44_5 ;
    input n5658;
    input n5657;
    input n5656;
    output \REG.mem_44_2 ;
    input n5655;
    input n5654;
    output \REG.mem_44_0 ;
    input n5653;
    output \REG.mem_43_15 ;
    input n5652;
    input n5651;
    output \REG.mem_43_13 ;
    input n5650;
    output \REG.mem_43_12 ;
    input n5649;
    output \REG.mem_43_11 ;
    input n5648;
    output \REG.mem_43_10 ;
    input n5647;
    output \REG.mem_43_9 ;
    input n5646;
    input n5645;
    output \REG.mem_43_7 ;
    input n5644;
    output \REG.mem_43_6 ;
    output \REG.mem_41_5 ;
    output \REG.mem_40_5 ;
    output \REG.mem_23_1 ;
    output \rd_addr_p1_w[0] ;
    output \REG.mem_35_11 ;
    input n5643;
    input n5642;
    input n5641;
    input n5640;
    output \REG.mem_43_2 ;
    input n5639;
    output \REG.mem_43_1 ;
    input n5638;
    input n5637;
    output \REG.mem_42_15 ;
    input n5636;
    input n5635;
    output \REG.mem_42_13 ;
    input n5634;
    output \REG.mem_42_12 ;
    input n5633;
    output \REG.mem_42_11 ;
    input n5632;
    output \REG.mem_42_10 ;
    input n5631;
    output \REG.mem_42_9 ;
    input n5630;
    input n5629;
    output \REG.mem_42_7 ;
    input n4916;
    output \REG.mem_31_6 ;
    output \REG.mem_23_2 ;
    output \REG.mem_38_11 ;
    output \REG.mem_39_11 ;
    output \REG.mem_37_11 ;
    output \REG.mem_36_11 ;
    input n5628;
    output \REG.mem_42_6 ;
    input n5627;
    input n5626;
    input n5625;
    input n5624;
    output \REG.mem_42_2 ;
    input n5623;
    output \REG.mem_42_1 ;
    input n5622;
    input n5621;
    output \REG.mem_41_15 ;
    input n5620;
    input n5619;
    output \REG.mem_41_13 ;
    input n5618;
    output \REG.mem_41_12 ;
    input n5617;
    output \REG.mem_41_11 ;
    input n5616;
    output \REG.mem_41_10 ;
    input n5615;
    output \REG.mem_41_9 ;
    input n5614;
    input n5613;
    output \REG.mem_41_7 ;
    output \REG.mem_3_2 ;
    input n5612;
    output \REG.mem_41_6 ;
    input n5611;
    input n5610;
    input n5609;
    input n5608;
    output \REG.mem_41_2 ;
    input n5607;
    output \REG.mem_41_1 ;
    input n5606;
    input n5605;
    output \REG.mem_40_15 ;
    input n5604;
    input n5603;
    output \REG.mem_40_13 ;
    input n5602;
    output \REG.mem_40_12 ;
    input n5601;
    output \REG.mem_40_11 ;
    input n5600;
    output \REG.mem_40_10 ;
    input n5599;
    output \REG.mem_40_9 ;
    input n5598;
    input n5597;
    output \REG.mem_40_7 ;
    output \REG.mem_25_9 ;
    input n4904;
    input n4903;
    input n4901;
    input n4899;
    input n5596;
    output \REG.mem_40_6 ;
    input n5595;
    input n5594;
    input n5593;
    input n5592;
    output \REG.mem_40_2 ;
    input n5591;
    output \REG.mem_40_1 ;
    input n5590;
    input n5589;
    input n5588;
    output \REG.mem_39_14 ;
    input n5587;
    input n5586;
    output \REG.mem_39_12 ;
    input n5585;
    input n5584;
    output \REG.mem_39_10 ;
    input n5583;
    output \REG.mem_39_9 ;
    input n5582;
    input n5581;
    input n4898;
    output \REG.mem_14_1 ;
    output \REG.mem_15_1 ;
    input DEBUG_5_c;
    output \REG.mem_13_1 ;
    output \REG.mem_12_1 ;
    output \REG.mem_3_3 ;
    input n5580;
    input n5579;
    input n5578;
    output \REG.mem_39_4 ;
    input n5577;
    input n5576;
    input n5575;
    output \REG.mem_39_1 ;
    input n5573;
    input n5572;
    input n5571;
    output \REG.mem_38_14 ;
    input n5570;
    input n5569;
    output \REG.mem_38_12 ;
    input n5568;
    input n5567;
    output \REG.mem_38_10 ;
    input n5566;
    output \REG.mem_38_9 ;
    input n5565;
    input n5564;
    input n5563;
    input n5562;
    input n5561;
    output \REG.mem_38_4 ;
    input n5560;
    input n5559;
    input n5558;
    output \REG.mem_38_1 ;
    input n5556;
    input n5555;
    input n5554;
    output \REG.mem_37_14 ;
    input n5553;
    input n5552;
    output \REG.mem_37_12 ;
    input n5551;
    input n5550;
    output \REG.mem_37_10 ;
    input n5549;
    output \REG.mem_37_9 ;
    output \REG.mem_25_13 ;
    output \REG.out_raw[15] ;
    output \REG.out_raw[14] ;
    output \REG.out_raw[13] ;
    output \REG.out_raw[12] ;
    output \REG.out_raw[11] ;
    input n5548;
    input n5547;
    input n5546;
    input n5545;
    input n5544;
    output \REG.mem_37_4 ;
    input n5543;
    input n5542;
    input n5541;
    output \REG.mem_37_1 ;
    input n5540;
    output \REG.out_raw[10] ;
    output \REG.out_raw[9] ;
    output \REG.out_raw[8] ;
    output \REG.out_raw[7] ;
    output \REG.out_raw[6] ;
    output \REG.out_raw[5] ;
    output \REG.out_raw[4] ;
    output \REG.out_raw[3] ;
    output \REG.out_raw[2] ;
    output \REG.out_raw[1] ;
    input n5526;
    input n5525;
    output \REG.mem_36_14 ;
    input n5524;
    input n5523;
    output \REG.mem_36_12 ;
    input n5522;
    input n5521;
    output \REG.mem_36_10 ;
    input n5520;
    output \REG.mem_36_9 ;
    input n5519;
    input n5518;
    input n5517;
    input n5516;
    output \rd_sig_diff0_w[2] ;
    input n5515;
    output \REG.mem_36_4 ;
    input n5514;
    input n5513;
    input n5512;
    output \REG.mem_36_1 ;
    input n5511;
    input n5507;
    input n5506;
    output \REG.mem_35_14 ;
    input n5505;
    input n5504;
    output \REG.mem_35_12 ;
    input n5503;
    input n5502;
    output \REG.mem_35_10 ;
    input n5501;
    output \REG.mem_35_9 ;
    input n5500;
    output \rd_sig_diff0_w[1] ;
    input n5499;
    output \REG.mem_35_7 ;
    input n5498;
    output \REG.mem_35_6 ;
    input n5497;
    output \REG.mem_35_5 ;
    input n5496;
    output \REG.mem_35_4 ;
    input n5495;
    input n5494;
    input n5493;
    output \REG.mem_35_1 ;
    input n5492;
    output \REG.mem_6_3 ;
    output \REG.mem_7_3 ;
    output \REG.mem_5_3 ;
    output \REG.mem_4_3 ;
    input n5441;
    input n5440;
    output \REG.mem_31_14 ;
    input n5439;
    input n5438;
    input n5437;
    output \REG.mem_25_1 ;
    input n5436;
    output \REG.mem_31_10 ;
    output n58;
    input n5435;
    output \REG.mem_31_9 ;
    input n5434;
    output \REG.mem_31_8 ;
    input n5433;
    input n5432;
    input n5431;
    input n5430;
    input n5429;
    input n5428;
    input n5427;
    output \REG.mem_31_1 ;
    input n5426;
    output n26;
    input DEBUG_1_c_c;
    output write_to_dc32_fifo_latched_N_425;
    input n5345;
    input n5344;
    output \REG.mem_25_14 ;
    input n5343;
    input n5342;
    input n5341;
    input n5340;
    output \REG.mem_25_10 ;
    input n5339;
    input n5338;
    output \REG.mem_25_8 ;
    input n5337;
    input n5336;
    input n5335;
    input n5334;
    input n5333;
    output \REG.mem_25_3 ;
    input n5332;
    input n5331;
    input n5330;
    output \REG.mem_25_0 ;
    output \REG.mem_14_15 ;
    output \REG.mem_15_15 ;
    output \REG.mem_6_13 ;
    output \REG.mem_7_13 ;
    input n5306;
    input n5305;
    output \REG.mem_23_14 ;
    input n5304;
    output \REG.mem_23_13 ;
    input n5303;
    input n5302;
    input n5301;
    output \REG.mem_23_10 ;
    input n5300;
    output \REG.mem_23_9 ;
    input n5299;
    input n5298;
    output \REG.mem_23_7 ;
    input n5297;
    output \REG.mem_23_6 ;
    input n5296;
    output \REG.mem_23_5 ;
    input n5295;
    output \REG.mem_23_4 ;
    input n5294;
    output \REG.mem_23_3 ;
    input n5293;
    input n5292;
    input n5290;
    output \REG.mem_23_0 ;
    output \rd_grey_sync_r[5] ;
    output \REG.mem_5_13 ;
    output \REG.mem_4_13 ;
    output \rd_grey_sync_r[4] ;
    output \rd_grey_sync_r[3] ;
    output \rd_grey_sync_r[2] ;
    output \rd_grey_sync_r[1] ;
    output \REG.mem_13_15 ;
    output \REG.mem_12_15 ;
    output n51;
    output n19;
    output \wr_addr_nxt_c[1] ;
    output \REG.mem_10_0 ;
    output \REG.mem_11_0 ;
    output \REG.mem_10_3 ;
    output \REG.mem_11_3 ;
    input n5224;
    input n5223;
    output \REG.mem_18_14 ;
    input n5222;
    output \REG.mem_18_13 ;
    input n5221;
    input n5220;
    output \REG.mem_9_3 ;
    output \REG.mem_8_3 ;
    output \REG.mem_9_0 ;
    output \REG.mem_8_0 ;
    output \REG.mem_10_13 ;
    output \REG.mem_11_13 ;
    output n52;
    output \REG.mem_9_13 ;
    output \REG.mem_8_13 ;
    output n20;
    input n5219;
    output \REG.mem_18_10 ;
    input n5218;
    output \REG.mem_18_9 ;
    input n5217;
    input n5216;
    input n5215;
    input n5214;
    output \REG.mem_18_5 ;
    input n5213;
    output \REG.mem_18_4 ;
    input n5212;
    output \REG.mem_18_3 ;
    input n5211;
    input n5210;
    input n5209;
    output \REG.mem_18_0 ;
    output \REG.mem_14_13 ;
    output \REG.mem_15_13 ;
    output \REG.mem_13_13 ;
    output \REG.mem_12_13 ;
    output \REG.mem_6_4 ;
    output \REG.mem_7_4 ;
    output \REG.mem_5_4 ;
    output \REG.mem_4_4 ;
    input get_next_word;
    input n5188;
    input n5186;
    output \REG.mem_16_14 ;
    input n5185;
    output \REG.mem_16_13 ;
    output \REG.mem_6_8 ;
    output \REG.mem_7_8 ;
    output \REG.mem_3_6 ;
    input n5184;
    output \REG.mem_5_8 ;
    output \REG.mem_4_8 ;
    output \REG.mem_6_2 ;
    output \REG.mem_7_2 ;
    output \REG.mem_5_2 ;
    output \REG.mem_4_2 ;
    output rd_fifo_en_w;
    input n5183;
    input n5182;
    output \REG.mem_16_10 ;
    input n5181;
    output \REG.mem_16_9 ;
    input n5180;
    input n5179;
    input n5178;
    input n5177;
    output \REG.mem_16_5 ;
    input n5176;
    output \REG.mem_16_4 ;
    output \REG.mem_3_12 ;
    input n5175;
    output \REG.mem_16_3 ;
    input n5174;
    input n5173;
    input n5172;
    output \REG.mem_16_0 ;
    input n5169;
    input n5168;
    input n5167;
    output n47;
    input n5166;
    output n15;
    input n5165;
    input n5164;
    output \REG.mem_15_10 ;
    input n5163;
    output \REG.mem_15_9 ;
    input n5162;
    input n5161;
    input n5160;
    output \REG.mem_15_6 ;
    input n5159;
    input n5158;
    input n5157;
    output \REG.mem_15_3 ;
    input n5156;
    output \REG.mem_15_2 ;
    input n5155;
    input n5154;
    output \REG.mem_15_0 ;
    input n5153;
    input n5152;
    output \REG.mem_6_6 ;
    output \REG.mem_7_6 ;
    input n5151;
    input n5150;
    input n5149;
    input n5148;
    output \REG.mem_14_10 ;
    input n5147;
    output \REG.mem_14_9 ;
    input n5146;
    input n5145;
    input n5144;
    output \REG.mem_14_6 ;
    output \REG.mem_4_6 ;
    output \REG.mem_5_6 ;
    input n5143;
    input n5142;
    input n5141;
    output \REG.mem_14_3 ;
    input n5140;
    output \REG.mem_14_2 ;
    input n5139;
    input n5138;
    output \REG.mem_14_0 ;
    input n5137;
    input n5136;
    input n5135;
    input n5134;
    input n5133;
    input n5132;
    output \REG.mem_13_10 ;
    output \REG.mem_13_9 ;
    output \REG.mem_12_9 ;
    input n5131;
    input n5130;
    input n5129;
    input n5128;
    output \REG.mem_13_6 ;
    input n5127;
    input n5126;
    input n5125;
    output \REG.mem_13_3 ;
    input n5124;
    output \REG.mem_13_2 ;
    input n5123;
    output \REG.mem_10_8 ;
    output \REG.mem_11_8 ;
    input n5122;
    output \REG.mem_13_0 ;
    input n5121;
    input n5120;
    input n5119;
    input n5118;
    output \REG.mem_3_9 ;
    output \REG.mem_9_8 ;
    output \REG.mem_8_8 ;
    input n5117;
    output \REG.mem_8_6 ;
    output \REG.mem_9_6 ;
    input n5116;
    output \REG.mem_12_10 ;
    output \REG.mem_10_6 ;
    output \REG.mem_11_6 ;
    output n53;
    output n21;
    input n5115;
    input n5114;
    input n5113;
    input n5112;
    output \REG.mem_12_6 ;
    output n50;
    input n5111;
    output n18;
    output \REG.mem_6_12 ;
    output \REG.mem_7_12 ;
    input n5110;
    input n5109;
    output \REG.mem_12_3 ;
    input n5108;
    output \REG.mem_12_2 ;
    output \REG.mem_4_12 ;
    output \REG.mem_5_12 ;
    output \REG.mem_10_2 ;
    output \REG.mem_11_2 ;
    input n5107;
    output \REG.mem_9_2 ;
    output \REG.mem_8_2 ;
    output n54;
    output n22;
    input n5106;
    output \REG.mem_12_0 ;
    output \rd_addr_nxt_c_6__N_498[3] ;
    input n5105;
    input n5104;
    input n5103;
    input n5102;
    output \REG.mem_11_12 ;
    input n5101;
    input n5100;
    output \REG.mem_11_10 ;
    input n5099;
    input n5098;
    input n5097;
    input n5096;
    input n5095;
    output \REG.mem_11_5 ;
    input n5094;
    input n5093;
    input n5092;
    input n5091;
    output \REG.mem_11_1 ;
    input n5090;
    input n5089;
    input n5088;
    output \rd_addr_nxt_c_6__N_498[5] ;
    input n5087;
    input n5086;
    output \REG.mem_10_12 ;
    input n5085;
    input n5084;
    output \REG.mem_10_10 ;
    input n5083;
    input n5082;
    input n5081;
    input n5080;
    input n5079;
    output \REG.mem_10_5 ;
    output \REG.mem_10_1 ;
    output \REG.mem_9_1 ;
    output \REG.mem_8_1 ;
    output \rd_addr_nxt_c_6__N_498[2] ;
    output n56;
    output n24;
    input n5078;
    output n55;
    output n23;
    input n5077;
    output n40;
    output n8;
    input n5076;
    input n5075;
    input n5074;
    input n5073;
    input n5072;
    input n5071;
    input n5070;
    output \REG.mem_9_12 ;
    input n5069;
    input n5068;
    output \REG.mem_9_10 ;
    input n5067;
    input n5066;
    input n5065;
    output n57;
    input n5064;
    output n25;
    input n5063;
    output \REG.mem_9_5 ;
    input n5062;
    input n5061;
    input n5060;
    input n5059;
    input n5057;
    input n5056;
    input n5055;
    input n5054;
    input n5053;
    output \REG.mem_8_12 ;
    input n5052;
    input n5051;
    output \REG.mem_8_10 ;
    input n5050;
    input n5049;
    input n5048;
    input n5047;
    input n5046;
    output \REG.mem_8_5 ;
    input n5045;
    input n5044;
    input n5043;
    input n5042;
    input n5041;
    input n5040;
    input n5039;
    input n5038;
    input n5037;
    input n5036;
    input n5035;
    output \REG.mem_7_10 ;
    input n5034;
    input n5033;
    input n5032;
    output \REG.mem_7_7 ;
    input n5031;
    input n5030;
    output \REG.mem_7_5 ;
    input n5029;
    input n5028;
    input n5027;
    input n5026;
    input n5025;
    output \REG.mem_7_0 ;
    input n5024;
    input n5023;
    input n5022;
    input n5021;
    input n5020;
    input n5019;
    output \REG.mem_6_10 ;
    input n5018;
    input n5017;
    input n5016;
    output \REG.mem_6_7 ;
    input n5015;
    input n5014;
    output \REG.mem_6_5 ;
    input n5013;
    input n5012;
    input n5011;
    input n5010;
    input n5009;
    output \REG.mem_6_0 ;
    input n5008;
    input n5007;
    input n5006;
    input n5005;
    input n5004;
    input n5003;
    output \REG.mem_5_10 ;
    input n5002;
    input n5001;
    input n5000;
    output \REG.mem_5_7 ;
    input n4999;
    input n4998;
    output \REG.mem_5_5 ;
    input n4997;
    input n4996;
    input n4995;
    input n4994;
    input n4993;
    output \REG.mem_5_0 ;
    input n4992;
    input n4991;
    input n4990;
    input n4989;
    input n4988;
    input n4987;
    output \REG.mem_4_10 ;
    input n4986;
    input n4985;
    input n4984;
    output \REG.mem_4_7 ;
    input n4983;
    input n4982;
    output \REG.mem_4_5 ;
    input n4981;
    input n4980;
    input n4979;
    input n4978;
    input n4977;
    output \REG.mem_4_0 ;
    input n4976;
    input n4975;
    input n4974;
    input n4973;
    input n4972;
    input n4971;
    output \REG.mem_3_10 ;
    input n4970;
    input n4969;
    output \REG.mem_3_8 ;
    output FT_OE_N_420;
    output n49;
    output n17;
    output n42;
    output n10;
    input n4968;
    output \REG.mem_3_7 ;
    input n4967;
    input n4966;
    output \REG.mem_3_5 ;
    input n4965;
    output n34;
    input n4964;
    input n4963;
    output n2;
    input n4962;
    input n4961;
    output \REG.mem_3_0 ;
    output n59;
    output n27;
    output n60;
    output n28;
    output n61;
    output n29;
    
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [6:0]rd_addr_r_c;   // src/fifo_dc_32_lut_gen.v(217[29:38])
    
    wire n12773, n13421, n11523, n11522, n13424, n43;
    wire [6:0]wr_addr_r;   // src/fifo_dc_32_lut_gen.v(196[29:38])
    
    wire \REG.mem_51_6 , n5778, \afull_flag_impl.af_flag_nxt_w , n12776, 
        \REG.mem_51_5 , n5777, \REG.mem_51_4 , n5776, \REG.mem_30_0 , 
        n12767, \REG.mem_29_0 , \REG.mem_28_0 , n12770, n13724, n13700, 
        n11022, \REG.mem_51_3 , n5775, \REG.mem_54_13 , n13415;
    wire [6:0]n1;
    
    wire n42_c, \REG.mem_34_2 , n5477, n11430, n11429, \REG.mem_17_8 , 
        n11393, \REG.mem_19_8 , n11394, \REG.mem_51_2 , n5774, \REG.mem_53_13 , 
        \REG.mem_52_13 , n13418, n11246, n11247, n12305, \REG.mem_2_13 , 
        n12425, \REG.mem_58_6 , \REG.mem_59_6 , n13409, n4950, \REG.mem_2_5 , 
        \REG.mem_56_6 , n11593, \REG.mem_51_1 , n5773, \REG.mem_62_11 , 
        n12761, \REG.mem_51_0 , n5772, \REG.mem_61_11 , \REG.mem_60_11 , 
        n11737, \REG.mem_34_1 , n5476, n12698, n13802;
    wire [31:0]\REG.out_raw_31__N_559 ;
    
    wire n12884, n13160, n13028, n13586, full_nxt_c_N_626, full_o, 
        n12992, n12824, n11391, n12962, n11392, n11531, n11532, 
        n13403, \REG.mem_34_0 , n12755, n13088, n13334, n11511, 
        n11510, n11595, n12788, n13286, n4949, \REG.mem_2_4 , n13082, 
        n13376, \REG.mem_33_0 , \REG.mem_32_0 , n11320, \REG.mem_54_10 , 
        n11520, n20_c, \REG.mem_52_10 , \REG.mem_53_10 , n11519, n4948, 
        \REG.mem_2_3 , \REG.mem_30_3 , n13397, n13484, n13748, n12800, 
        n13238, n11116, n12638, n11184, \REG.mem_29_3 , \REG.mem_28_3 , 
        n11077, n12842, n12734, n13532, \REG.mem_49_7 , n11474, 
        \REG.mem_51_7 , n11475, \REG.mem_54_7 , n11505, n4947, \REG.mem_2_2 , 
        \REG.mem_52_7 , \REG.mem_53_7 , n11504, n11068, n12749, n5474, 
        \REG.mem_1_13 , \REG.mem_0_13 , n11815, n11065, n11059, n11137, 
        n11555, n11556, n13391, \REG.mem_49_10 , n11516, \REG.mem_51_10 , 
        n11517, n11870, n11871, n12743, n11541, n11540, n13394;
    wire [6:0]wr_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(200[30:42])
    
    wire wr_sig_mv_w;
    wire [6:0]wr_grey_w;   // src/fifo_dc_32_lut_gen.v(203[38:47])
    
    wire n11868, n11867, n12746, \REG.mem_22_8 , n11442, \REG.mem_58_9 , 
        \REG.mem_59_9 , n12419, \REG.mem_20_8 , \REG.mem_21_8 , n11441, 
        \REG.mem_26_5 , \REG.mem_27_5 , n13385, n5672, \REG.mem_24_5 , 
        n13388;
    wire [6:0]rd_grey_w;   // src/fifo_dc_32_lut_gen.v(224[38:47])
    
    wire \REG.mem_26_15 , \REG.mem_27_15 , n12737, \REG.mem_24_15 , 
        n12740, n12326, n13850, n11568, n4946, \REG.mem_2_1 , n12542, 
        n12362, n11567, n13379, n12650, n11016, n12731, empty_nxt_c_N_629, 
        n13382, n4945, \REG.mem_2_0 , n4944, \REG.mem_0_0 , n13070, 
        n11586, n13373, n4943, \REG.mem_0_1 , n13154, n12656, n11553, 
        n11952, n11951, n11562, n13052, n13367, n11623, n11632, 
        n12725, n11230, \REG.mem_56_9 , n12422, n11611, n11608, 
        n11743, n13778, n13754, n11019, n11894, n11895, n12719, 
        \REG.mem_34_3 , n13361, \REG.mem_33_3 , \REG.mem_32_3 , n11080, 
        n11883, n11882, n12722, n13355, n13358, \REG.mem_24_2 , 
        n11885, n11864, n11865, n12713, n39, \REG.mem_17_15 , n5208, 
        \REG.mem_17_14 , n5207, \REG.mem_26_2 , \REG.mem_27_2 , n11886, 
        \REG.mem_17_13 , n5206, \REG.mem_2_11 , n13349, n4941, \REG.mem_0_2 , 
        \REG.mem_1_11 , \REG.mem_0_11 , n11856, n11855, n12716, \REG.mem_30_2 , 
        n11898, \REG.mem_28_2 , \REG.mem_29_2 , n11897, \REG.mem_51_12 , 
        n12707, \REG.mem_17_12 , n5205, n13343, \REG.mem_17_11 , n5204, 
        n11232, n11231, n12308, \REG.mem_49_12 , n12710, n11965, 
        n11971, n12311, n12299, n12701, n11858, \REG.mem_17_10 , 
        n5203, n11859, \REG.mem_62_6 , n13337, n4940, \REG.mem_0_3 , 
        n12704, n11862, n11012, n12470, n12695, \REG.mem_17_9 , 
        n5202, n5201, n12413, \REG.mem_17_7 , n5200, n11010, n11009, 
        n11861, n11852, n11853, n12689, \REG.mem_61_6 , \REG.mem_60_6 , 
        n11614, \REG.mem_17_6 , n5199, n11850, n11849, n12692, \REG.mem_17_5 , 
        n5198, \REG.mem_17_4 , n5197, n13076, n13331, n11583, n13064, 
        \REG.mem_17_3 , n5196, n12683, \REG.mem_17_2 , n5195, \REG.mem_17_1 , 
        n5194, n11171, n11172, n13325, n11169, n11168, n11250, 
        n12686, \REG.mem_17_0 , n5193, n11948, n11949, n12677, \REG.mem_19_12 , 
        n13319, \REG.mem_1_1 , n12416, \REG.mem_19_15 , n5240, n13322, 
        \REG.mem_19_14 , n5239, \REG.mem_19_13 , n5238, n11943, n11942, 
        n12680, n5237, \REG.mem_19_11 , n5236, \REG.mem_19_10 , n5235, 
        \REG.mem_19_9 , n5234, n5233, n11909, n11910, n12671, n11198, 
        n11199, n13313, \REG.mem_19_7 , n5232, n11907, n11906, n12674, 
        \REG.mem_19_6 , n5231, \REG.mem_30_15 , n12665, n11193, n11192, 
        n11256, \REG.mem_19_5 , n5230, \REG.mem_19_4 , n5229, \REG.mem_19_3 , 
        n5228, \REG.mem_29_15 , \REG.mem_28_15 , n12668, n13307, n11086, 
        n11656, n11668, n12659, n11653, n11644, n11755, \REG.mem_19_2 , 
        n5227, n13301, \REG.mem_19_1 , n5226, n12653, n11089, n11714, 
        n11715, n12647, \REG.mem_19_0 , n5225, n11694, n11693, \REG.mem_58_0 , 
        \REG.mem_59_0 , n13295, \REG.mem_56_0 , n13298, n11681, n11682, 
        n12641, n13289, n11637, n11636, n12644, \REG.mem_62_12 , 
        n12407, n45, \REG.mem_20_15 , n5256, \REG.mem_20_14 , n5255, 
        \REG.mem_20_13 , n5254, \REG.mem_20_12 , n5253, \REG.mem_20_11 , 
        n5252, \REG.mem_20_10 , n5251, n10993, n10996, n12635, n11049, 
        n13283, n12016, n12010, \REG.mem_20_9 , n5250, \REG.mem_54_12 , 
        n12629, n11004, \REG.mem_53_12 , \REG.mem_52_12 , n12632, 
        n11219, n11220, n13277, \REG.mem_34_15 , n12623, \REG.mem_33_15 , 
        \REG.mem_32_15 , n12626, n11217, n11216, n11259, \REG.mem_2_15 , 
        n13271, n5249, \REG.mem_20_7 , n5248, \REG.mem_1_15 , \REG.mem_0_15 , 
        n13274, n4935, \REG.mem_0_4 , \REG.mem_51_9 , n12617, n4934, 
        \REG.mem_0_5 , \REG.mem_49_9 , n12620, \REG.mem_20_6 , n5247, 
        \REG.mem_20_5 , n5246, \REG.mem_1_4 , n12302, n12293, \REG.mem_20_4 , 
        n5245, \REG.mem_20_3 , n5244, n13265, n12296, n12335, n12338, 
        n12329, n11692, n11701, n12611, n11104, \REG.mem_20_2 , 
        n5243, \REG.mem_20_1 , n5242, n12323, \REG.mem_24_7 , \REG.mem_22_12 , 
        n13259, \REG.mem_20_0 , n5241, n11677, n11674, n11764, n11158, 
        n11176, n12317, n47_c, \REG.mem_21_15 , n5273, \REG.mem_21_12 , 
        n13262, \REG.mem_61_12 , \REG.mem_60_12 , n12410, n11959, 
        n12314, \REG.mem_21_14 , n5272, \REG.mem_21_13 , n5271, n5270, 
        \REG.mem_21_11 , n5269, \REG.mem_21_10 , n5268, \REG.mem_21_9 , 
        n5267, n12605, n11455, n11488, n12287, \REG.mem_30_13 , 
        n13253, n11332, \REG.mem_29_13 , \REG.mem_28_13 , n13256, 
        n5266, n11722, n12599, n13247, n11110, \REG.mem_21_7 , n5265, 
        \REG.mem_21_6 , n5264, \REG.mem_21_5 , n5263, \REG.mem_21_4 , 
        n5262, \REG.mem_21_3 , n5261, n13241, n11719, n11710, n11767, 
        \REG.mem_49_3 , n11113, \REG.mem_21_2 , n5260, \REG.mem_21_1 , 
        n5259, n12593, \REG.mem_21_0 , n5257, n49_c, \REG.mem_22_15 , 
        n5289, \REG.mem_22_14 , n5288, \REG.mem_22_13 , n5287, n11996, 
        n11997, n13235, n11335, n11991, n11990, n5286, \REG.mem_22_11 , 
        n5285, \REG.mem_22_10 , n5284, \REG.mem_22_9 , n5283, n5282, 
        \REG.mem_22_7 , n5281, \REG.mem_22_6 , n5280, \REG.mem_22_5 , 
        n5279, \REG.mem_22_4 , n5278, \REG.mem_22_3 , n5277, \REG.mem_22_2 , 
        n5276, n13229, \REG.mem_22_1 , n5275, \REG.mem_22_0 , n5274, 
        n53_c, n5329, n11728, n11785, n12401, \REG.mem_24_14 , n5328, 
        \REG.mem_24_13 , n5327, n11704, n11659, \REG.mem_24_12 , n5326, 
        \REG.mem_58_13 , \REG.mem_59_13 , n13223, \REG.mem_24_11 , n5325, 
        n12581, n12584, \REG.mem_56_13 , n13226, n11240, n11241, 
        n13217, \REG.mem_24_10 , n5324, n4933, \REG.mem_0_6 , \REG.mem_24_9 , 
        n5323, n11238, n11237, n11262, \REG.mem_24_8 , n5322, n5321, 
        n13211, n12575, \REG.mem_24_6 , n5320, \REG.mem_49_1 , n13214, 
        n13205, \REG.mem_49_15 , n5752, n12956, n11383, \REG.mem_49_14 , 
        n5751, n5319, \REG.mem_24_4 , n5318, \REG.mem_24_3 , n5317, 
        n5316, n11143, \REG.mem_24_1 , n5315, \REG.mem_24_0 , n5307, 
        \REG.mem_49_13 , n5750, n57_c, n5361, n5749, \REG.mem_26_14 , 
        n5360, \REG.mem_49_11 , n5748, \REG.mem_30_5 , n13199, n5747, 
        \REG.mem_29_5 , \REG.mem_28_5 , n13202, n5746, \REG.mem_49_8 , 
        n5745, \REG.mem_26_12 , \REG.mem_27_12 , n13193, \REG.mem_26_13 , 
        n5359, n5358, n5744, n13196, n12395, \REG.mem_49_6 , n5743, 
        \REG.mem_49_5 , n5742, \REG.mem_26_11 , n5357, \REG.mem_49_4 , 
        n5741, n4932, \REG.mem_0_7 , n5740;
    wire [6:0]wp_sync2_r;   // src/fifo_dc_32_lut_gen.v(223[37:47])
    wire [6:0]wp_sync_w;   // src/fifo_dc_32_lut_gen.v(226[30:39])
    
    wire \REG.mem_26_10 , n5356, \REG.mem_26_9 , n5355, \REG.mem_26_8 , 
        n5354, \REG.mem_26_7 , n5353, \REG.mem_49_2 , n5739, \REG.mem_26_6 , 
        n5352, n13187, n5738, n5351, n6044, n6042, n13190, \REG.mem_49_0 , 
        n5737, \REG.mem_34_13 , n13181, n11947, n12551, n4931, \REG.mem_0_8 , 
        n12554, \REG.mem_33_13 , \REG.mem_32_13 , n13184, \REG.mem_27_6 , 
        n13175, \REG.mem_26_4 , n5350, n12545, \REG.mem_26_3 , n5349, 
        n6005, \REG.mem_62_15 , n6004, \REG.mem_62_14 , n6003, \REG.mem_62_13 , 
        n6002, n4930, \REG.mem_0_9 , n11272, n12398, n11146, n5348, 
        \REG.mem_56_4 , n12539, \REG.mem_58_4 , \REG.mem_59_4 , n12533, 
        n4929, \REG.mem_0_10 , n4928, n11545, n11530, n6001, n6000, 
        \REG.mem_62_10 , n5999, \REG.mem_62_9 , n5998, \REG.mem_62_8 , 
        n5997, \REG.mem_62_7 , n5996, n5995, \REG.mem_62_5 , n5994, 
        \REG.mem_62_4 , n5993, \REG.mem_62_3 , n5992, \REG.mem_62_2 , 
        n5991, \REG.mem_62_1 , n5990, \REG.mem_62_0 , n5986, \REG.mem_61_15 , 
        n5985, \REG.mem_61_14 , \REG.mem_26_1 , n5347, n12527, n13169, 
        n12530, \REG.mem_26_0 , n5346, n11125, n11128, n12521, n11119, 
        n11149, n12515, n11131, n5984, \REG.mem_61_13 , n5983, n5982, 
        n5981, \REG.mem_61_10 , n5980, \REG.mem_61_9 , n5979, \REG.mem_61_8 , 
        n5978, \REG.mem_61_7 , n5977, n5976, \REG.mem_61_5 , n5975, 
        \REG.mem_61_4 , n5974, \REG.mem_61_3 , n5973, \REG.mem_61_2 , 
        n5972, \REG.mem_61_1 , n5971, \REG.mem_61_0 , n5969, \REG.mem_60_15 , 
        \REG.mem_27_11 , n13163, n59_c, n5377, \REG.mem_27_14 , n5376, 
        \REG.mem_58_12 , \REG.mem_59_12 , n12509, \REG.mem_60_4 , n12878, 
        n13157, \REG.mem_56_12 , n12512, \REG.mem_27_13 , n5375, n13142, 
        n13148, n12872, n5968, \REG.mem_60_14 , n5967, \REG.mem_60_13 , 
        n5966, n5965, n5964, \REG.mem_60_10 , n5963, \REG.mem_60_9 , 
        n5962, \REG.mem_60_8 , n5961, \REG.mem_60_7 , n5960, n5959, 
        \REG.mem_60_5 , n5958, n5957, \REG.mem_60_3 , n5956, \REG.mem_60_2 , 
        n5955, \REG.mem_60_1 , n5954, \REG.mem_60_0 ;
    wire [6:0]rp_sync2_r;   // src/fifo_dc_32_lut_gen.v(202[37:47])
    
    wire n5944, \REG.mem_59_15 , n5943, \REG.mem_59_14 , n5942, n5941, 
        n5940, \REG.mem_59_11 , n5939, \REG.mem_59_10 , n5938, n5937, 
        \REG.mem_59_8 , \REG.mem_54_9 , n12503, n5374, \REG.mem_53_9 , 
        \REG.mem_52_9 , n12506, n5936, \REG.mem_59_7 , n5935, n13151, 
        n5934, \REG.mem_59_5 , n5933, n5932, \REG.mem_59_3 , n5931, 
        \REG.mem_59_2 , n5930, \REG.mem_59_1 , n5929, n5925, n5922, 
        n5920, n5919, \REG.mem_58_15 , n5918, \REG.mem_58_14 , n4927, 
        \REG.mem_0_12 , n12497, n11093, n11094, n13145, n5373, n5917, 
        n5916, n5915, \REG.mem_58_11 , n5914, \REG.mem_58_10 , n5913, 
        n5912, \REG.mem_58_8 , n5911, \REG.mem_58_7 , n5910, n5909, 
        \REG.mem_58_5 , n5908, n5907, \REG.mem_58_3 , n5906, \REG.mem_58_2 , 
        n5905, \REG.mem_58_1 , n5904, n11001, n11000, \REG.mem_27_10 , 
        n5372, n13859, n11389, \REG.mem_27_9 , n5371, n12023, n12024, 
        n13139, \REG.mem_27_8 , n5370, n5884, \REG.mem_56_15 , n5883, 
        \REG.mem_56_14 , n5882, n5881, n5880, \REG.mem_56_11 , n5879, 
        \REG.mem_56_10 , n5878, n5877, \REG.mem_56_8 , n5876, \REG.mem_56_7 , 
        n5875, n5874, \REG.mem_56_5 , n5873, n5872, \REG.mem_56_3 , 
        n5871, \REG.mem_56_2 , n5870, \REG.mem_56_1 , \REG.mem_32_8 , 
        \REG.mem_33_8 , \REG.mem_34_8 , n12012, n12011, n13853, n5865, 
        n10137, n10138, n10136, n10135, n10090, n10091, n10134, 
        n10133;
    wire [6:0]rd_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(221[30:42])
    
    wire n10144, n10143;
    wire [6:0]n1_adj_45;
    
    wire n10101, n10979, n5835, \REG.mem_54_15 , n5834, \REG.mem_54_14 , 
        n5833, n5832, n5831, \REG.mem_54_11 , n5830, n5829, n5828, 
        \REG.mem_54_8 , n5827, n5826, \REG.mem_54_6 , n5825, \REG.mem_54_5 , 
        n5824, \REG.mem_54_4 , n5823, \REG.mem_54_3 , n5822, \REG.mem_54_2 , 
        n5821, \REG.mem_54_1 ;
    wire [6:0]rp_sync_w;   // src/fifo_dc_32_lut_gen.v(205[30:39])
    
    wire n10100, n10951, n10142, n10925, n10099, n2_adj_22;
    wire [6:0]wr_sig_diff0_w;   // src/fifo_dc_32_lut_gen.v(212[30:44])
    
    wire n10098, \REG.mem_27_4 , \REG.mem_32_2 , \REG.mem_33_2 , \REG.mem_30_4 , 
        n5820, \REG.mem_54_0 , n5819, \REG.mem_53_15 , n5818, \REG.mem_53_14 , 
        n5817, n5816, n5815, \REG.mem_53_11 , n5814, n5813, n5812, 
        \REG.mem_53_8 , n5811, n5810, \REG.mem_53_6 , n5809, \REG.mem_53_5 , 
        n5808, \REG.mem_53_4 , n5807, \REG.mem_53_3 , n5806, \REG.mem_53_2 , 
        n5805, \REG.mem_53_1 , \REG.mem_28_4 , \REG.mem_29_4 , n10141, 
        n5804, \REG.mem_53_0 , n5803, \REG.mem_52_15 , n5802, \REG.mem_52_14 , 
        n5801, n5800, n5799, \REG.mem_52_11 , n5798, n5797, n5796, 
        \REG.mem_52_8 , n5795, n5794, \REG.mem_52_6 , n5793, \REG.mem_52_5 , 
        n5792, \REG.mem_52_4 , n5791, \REG.mem_52_3 , n5790, \REG.mem_52_2 , 
        n5789, \REG.mem_52_1 , n13133, \REG.mem_27_7 , n5369, n10097, 
        n5788, \REG.mem_52_0 , n5787, \REG.mem_51_15 , n5786, \REG.mem_51_14 , 
        n5785, \REG.mem_51_13 , n5784, n5783, \REG.mem_51_11 , n5782, 
        n5781, n5780, \REG.mem_51_8 , n5779, n10096, n10140, n10095;
    wire [6:0]rd_sig_diff0_w;   // src/fifo_dc_32_lut_gen.v(233[30:44])
    
    wire n10094, \REG.mem_0_14 , \REG.mem_1_14 , \REG.mem_2_14 , n10139, 
        n12446, n12386, n10093, n13136, \REG.mem_30_7 , n13847, 
        \REG.mem_29_7 , \REG.mem_28_7 , n4926, n4925, n12368, n12350, 
        n12479, n4924, n12482, n12380, n13841, \REG.mem_30_12 , 
        n13127, n13814, n11401, n5368, \REG.mem_29_12 , \REG.mem_28_12 , 
        n13130, n13121, n13835, n11025, n13829, n5367, n5366, 
        n12467, n11407, \REG.mem_30_11 , n13115, \REG.mem_29_11 , 
        \REG.mem_28_11 , n12461, n13823, n13109, \REG.mem_27_3 , n5365, 
        n13112, n5364, \REG.mem_27_1 , n5363, \REG.mem_27_0 , n5362, 
        n12464, n12320, n61_c, n5393, \REG.mem_28_14 , n5392, n5391, 
        n10092, n13817, n5390, n11419, \REG.mem_34_11 , n13103, 
        \REG.mem_33_11 , \REG.mem_32_11 , \genblk16.rd_prev_r , n5389, 
        n12389, n11302, n12434, n12455, n12458, \REG.mem_30_6 , 
        n12449, n13811, \REG.mem_29_6 , \REG.mem_28_6 , n12452, n13097, 
        n4915, n4914, \REG.mem_1_6 , \REG.mem_28_10 , n5388, \REG.mem_28_9 , 
        n5387, n12830, n13091, n12443, \REG.mem_1_2 , n4912, \REG.mem_1_12 , 
        n12854, n12914, n13094, n13805, \REG.mem_28_8 , n5386, n4905, 
        \REG.mem_1_7 , n5385, n4902, n4900, \REG.mem_1_8 , n13085, 
        n13799, n6_adj_23, n12431, n13040, n13793, \REG.mem_1_3 , 
        n11035, n10254, n13046, n11559, n13079, n11550, n13034, 
        n5384, n5383, n5382, n5381, n5380, \REG.mem_28_1 , n5379, 
        n5378, n63, n5409, \REG.mem_29_14 , n5408, n12392, n5407, 
        n5406, n5405, \REG.mem_29_10 , n5404, n12341, n13787, n11440, 
        \REG.mem_29_9 , n5403, n13073, n13781, \REG.mem_29_8 , n5402, 
        n13784, n5401, n13067, n5400, n13775, n5399, n5398, n5397, 
        n5396, n5490, n5489, \REG.mem_34_14 , n5488, n5487, \REG.mem_34_12 , 
        n5486, n5485, \REG.mem_34_10 , n5484, \REG.mem_34_9 , \REG.mem_29_1 , 
        n5395, n5394, n65, n5425, \REG.mem_30_14 , n5424, n5423, 
        n5422, n5421, n13769, n5483, n5482, \REG.mem_34_7 , n5481, 
        \REG.mem_34_6 , n5480, \REG.mem_34_5 , n5479, \REG.mem_34_4 , 
        n5478, n5473, n5472, \REG.mem_33_14 , n5471, n5470, \REG.mem_33_12 , 
        n5469, n5468, \REG.mem_33_10 , \REG.mem_30_10 , n5420, n12020, 
        \REG.mem_30_9 , n5419, n13061, \REG.mem_30_8 , n5418, n13763, 
        n11041, n5467, \REG.mem_33_9 , n5466, n5465, \REG.mem_33_7 , 
        n5464, \REG.mem_33_6 , n5463, \REG.mem_33_5 , n5462, \REG.mem_33_4 , 
        n5461, n5460, n5459, \REG.mem_33_1 , n5458, n5457, n5456, 
        \REG.mem_32_14 , n5455, n5454, \REG.mem_32_12 , n5453, n11412, 
        n11411, n5417, n11285, n11286, n13055, n5452, \REG.mem_32_10 , 
        n5416, n5451, \REG.mem_32_9 , n5450, n5449, \REG.mem_32_7 , 
        n5448, \REG.mem_32_6 , n5447, \REG.mem_32_5 , n5446, \REG.mem_32_4 , 
        n5445, n5444, n5443, \REG.mem_32_1 , n5442, n13757, n11283, 
        n11282, n13058, n5415, n5414, n36, n11489, n11490, n13049, 
        n5413, n5412, n11478, n11477, \REG.mem_30_1 , n5411, n13751, 
        n11450, n11451, n13043, n5410, n11448, n11447, n38, n11243, 
        n11244, n13037, n11921, n11922, n13745, n11901, n11900, 
        n11202, n11201, n13739, n11464, n12938, n12812, n13733, 
        n4884, \REG.mem_1_0 , n11423, n11424, n13031, n11941, n11415, 
        n11414, n13727, n13010, n11472, n13025, n12344, n13721, 
        n11460, n12986, n11402, n11403, n13019, n11385, n11384, 
        n13022, n13013, n13715, n13016, n11905, n13709, n12290, 
        n17_c, n11204, n11205, n13007, n13703, n11482, n11163, 
        n11162, n13697, n13691, n13001, n11485, n13004, n40_c, 
        n12995, n13685, n11044, n12998, n13679, n15_c, n4274, 
        n10889, n10899, n13673, n11968, n4298, n10_c, n13667, 
        n8_adj_25, n12, n10887, n10985, n4960, n12989, n13661, 
        n13664, n11072, n11073, n12983, n10258, n4959, n4958, 
        \REG.mem_2_12 , n4957, n13655, \REG.mem_2_6 , n4956, n13658, 
        \REG.mem_2_10 , n4955, n12383, \REG.mem_2_9 , n4954, n11936, 
        n11937, n13649, n12377, \REG.mem_2_8 , n4953, \REG.mem_2_7 , 
        n4952, n11037, n11036, n11874, n11873, n4951;
    wire [6:0]rd_addr_nxt_c_6__N_498;
    
    wire n13643, n4879, n13637, n11500, n18_c, n12977, n11927, 
        n11928, n13631, n11919, n11918, n11052, \REG.mem_1_10 , 
        n4831, n12971, n13625, n12974, n13619, n12965, n11279, 
        n11280, n12959, \REG.mem_1_9 , n4833, n13622, n4867, n11253, 
        n11252, n4832, n13613, n11977, n11210, n11211, n12953, 
        n11187, n11186, n13607, n11983, \REG.mem_1_5 , n4835, n4837, 
        n13601, n4861, n12371, n4868, n12947, n13604, n11122, 
        n12941, n11197, n13, n11432, n11433, n13595, n12374, n12935, 
        n14, n11421, n11420, n11514, n13589, n11989, n35, n12929, 
        n12365, n12923, n12926, n13583, n4866, n12917, n11493, 
        n11492, n13577, n12920, n12911, n12905, n13571, n12899, 
        n12836, n13565, n11995, n23_c, n12893, n13559, n11575, 
        n13553, n12887, n11056, n12890, n12_adj_33, n13547, n12359, 
        n11914, n12866, n12881, n11249, n13541, n11234, n11235, 
        n12875, n13535, n11226, n11225, n11, n11213, n11214, n12869, 
        n13529, n11208, n11207, n11189, n11190, n12863, n11178, 
        n11177, n11028, n11027, n12353, n12857, n11435, n11436, 
        n13523, n11427, n11426, n13517, n13511, n12851, n13505, 
        n12356, n11468, n11469, n13499, n10845, n11457, n11456, 
        full_max_w, n12845, n10849, n10881, n12_adj_35, n3_adj_36, 
        n6_adj_37, n10947, n12032, n12033, n11507, n11508, n13493, 
        n11496, n11495, n13487, n13490, n11070, n12839, n11888, 
        n11889, n13481, n11877, n12833, n13475, n9, n12827, n13469, 
        n12821, n13472, n12815, n11915, n11916, n13463, n11892, 
        n11891, n12347, n12809, n13457, n13460, n12026, n12027, 
        n13451, n11984, n11985, n12797, n11973, n11972, n13454, 
        n11979, n11978, n13445, n13448, n12791, n13439, n12021, 
        n12785, n13442, n12003, n12002, n12779, n11465, n11466, 
        n13433, n12782, n11445, n11444, n11537, n11538, n13427, 
        n11535, n11534, n11546, n11547, n11904, n11574, n11913;
    
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10856 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_5 ), 
            .I2(\REG.mem_15_5 ), .I3(rd_addr_r_c[1]), .O(n12773));
    defparam rd_addr_r_0__bdd_4_lut_10856.LUT_INIT = 16'he4aa;
    SB_LUT4 n13421_bdd_4_lut (.I0(n13421), .I1(n11523), .I2(n11522), .I3(rd_addr_r_c[2]), 
            .O(n13424));
    defparam n13421_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4395_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_51_6 ), .O(n5778));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4395_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFSR \afull_flag_impl.af_flag_ext_r_121  (.Q(dc32_fifo_almost_full), 
            .C(FIFO_CLK_c), .D(\afull_flag_impl.af_flag_nxt_w ), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(410[29] 422[32])
    SB_LUT4 n12773_bdd_4_lut (.I0(n12773), .I1(\REG.mem_13_5 ), .I2(\REG.mem_12_5 ), 
            .I3(rd_addr_r_c[1]), .O(n12776));
    defparam n12773_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4394_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_51_5 ), .O(n5777));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4394_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4393_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_51_4 ), .O(n5776));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4393_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10851 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_0 ), 
            .I2(\REG.mem_31_0 ), .I3(rd_addr_r_c[1]), .O(n12767));
    defparam rd_addr_r_0__bdd_4_lut_10851.LUT_INIT = 16'he4aa;
    SB_LUT4 n12767_bdd_4_lut (.I0(n12767), .I1(\REG.mem_29_0 ), .I2(\REG.mem_28_0 ), 
            .I3(rd_addr_r_c[1]), .O(n12770));
    defparam n12767_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9184_3_lut (.I0(n13724), .I1(n13700), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11022));
    defparam i9184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4392_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_51_3 ), .O(n5775));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4392_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11405 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_13 ), 
            .I2(\REG.mem_55_13 ), .I3(rd_addr_r_c[1]), .O(n13415));
    defparam rd_addr_r_0__bdd_4_lut_11405.LUT_INIT = 16'he4aa;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i3_1_lut (.I0(rd_addr_r_c[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4094_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_34_2 ), .O(n5477));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4094_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9592_3_lut (.I0(\REG.mem_38_7 ), .I1(\REG.mem_39_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11430));
    defparam i9592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9591_3_lut (.I0(\REG.mem_36_7 ), .I1(\REG.mem_37_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11429));
    defparam i9591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9555_3_lut (.I0(\REG.mem_16_8 ), .I1(\REG.mem_17_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11393));
    defparam i9555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9556_3_lut (.I0(\REG.mem_18_8 ), .I1(\REG.mem_19_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11394));
    defparam i9556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4391_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_51_2 ), .O(n5774));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4391_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13415_bdd_4_lut (.I0(n13415), .I1(\REG.mem_53_13 ), .I2(\REG.mem_52_13 ), 
            .I3(rd_addr_r_c[1]), .O(n13418));
    defparam n13415_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10597 (.I0(rd_addr_r_c[1]), .I1(n11246), 
            .I2(n11247), .I3(rd_addr_r_c[2]), .O(n12305));
    defparam rd_addr_r_1__bdd_4_lut_10597.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10568 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_13 ), 
            .I2(\REG.mem_3_13 ), .I3(rd_addr_r_c[1]), .O(n12425));
    defparam rd_addr_r_0__bdd_4_lut_10568.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11385 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_6 ), 
            .I2(\REG.mem_59_6 ), .I3(rd_addr_r_c[1]), .O(n13409));
    defparam rd_addr_r_0__bdd_4_lut_11385.LUT_INIT = 16'he4aa;
    SB_DFF i245_246 (.Q(\REG.mem_2_5 ), .C(FIFO_CLK_c), .D(n4950));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13409_bdd_4_lut (.I0(n13409), .I1(\REG.mem_57_6 ), .I2(\REG.mem_56_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11593));
    defparam n13409_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4390_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_51_1 ), .O(n5773));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4390_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10846 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_11 ), 
            .I2(\REG.mem_63_11 ), .I3(rd_addr_r_c[1]), .O(n12761));
    defparam rd_addr_r_0__bdd_4_lut_10846.LUT_INIT = 16'he4aa;
    SB_LUT4 i4389_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_51_0 ), .O(n5772));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4389_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12761_bdd_4_lut (.I0(n12761), .I1(\REG.mem_61_11 ), .I2(\REG.mem_60_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11737));
    defparam n12761_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4093_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_34_1 ), .O(n5476));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4093_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9194_3_lut (.I0(n12698), .I1(n13802), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [2]));
    defparam i9194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9437_3_lut (.I0(n12884), .I1(n13160), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [4]));
    defparam i9437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9689_3_lut (.I0(n13028), .I1(n13586), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [5]));
    defparam i9689_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR full_ext_r_117 (.Q(full_o), .C(FIFO_CLK_c), .D(full_nxt_c_N_626), 
            .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 i9553_3_lut (.I0(n12992), .I1(n12824), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11391));
    defparam i9553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9554_3_lut (.I0(n12962), .I1(n11391), .I2(rd_addr_r_c[3]), 
            .I3(GND_net), .O(n11392));
    defparam i9554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11390 (.I0(rd_addr_r_c[1]), .I1(n11531), 
            .I2(n11532), .I3(rd_addr_r_c[2]), .O(n13403));
    defparam rd_addr_r_1__bdd_4_lut_11390.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10841 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_0 ), 
            .I2(\REG.mem_35_0 ), .I3(rd_addr_r_c[1]), .O(n12755));
    defparam rd_addr_r_0__bdd_4_lut_10841.LUT_INIT = 16'he4aa;
    SB_DFFE \REG.out_raw__i1  (.Q(\REG.out_raw[0] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [0]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_LUT4 i9779_3_lut (.I0(n13088), .I1(n13334), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [7]));
    defparam i9779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13403_bdd_4_lut (.I0(n13403), .I1(n11511), .I2(n11510), .I3(rd_addr_r_c[2]), 
            .O(n11595));
    defparam n13403_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9260_3_lut (.I0(n12788), .I1(n13286), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [8]));
    defparam i9260_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i242_243 (.Q(\REG.mem_2_4 ), .C(FIFO_CLK_c), .D(n4949));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9764_3_lut (.I0(n13082), .I1(n13376), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [10]));
    defparam i9764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12755_bdd_4_lut (.I0(n12755), .I1(\REG.mem_33_0 ), .I2(\REG.mem_32_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11320));
    defparam n12755_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9682_3_lut (.I0(\REG.mem_54_10 ), .I1(\REG.mem_55_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11520));
    defparam i9682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i76_2_lut_3_lut_4_lut (.I0(n20_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n62));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i76_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i9681_3_lut (.I0(\REG.mem_52_10 ), .I1(\REG.mem_53_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11519));
    defparam i9681_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i239_240 (.Q(\REG.mem_2_3 ), .C(FIFO_CLK_c), .D(n4948));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i75_2_lut_3_lut_4_lut (.I0(n20_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n30));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i75_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11380 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_3 ), 
            .I2(\REG.mem_31_3 ), .I3(rd_addr_r_c[1]), .O(n13397));
    defparam rd_addr_r_0__bdd_4_lut_11380.LUT_INIT = 16'he4aa;
    SB_LUT4 i10097_3_lut (.I0(n13484), .I1(n13748), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [12]));
    defparam i10097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9278_3_lut (.I0(n12800), .I1(n13238), .I2(rd_addr_r_c[3]), 
            .I3(GND_net), .O(n11116));
    defparam i9278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9346_3_lut (.I0(n11116), .I1(n12638), .I2(rd_addr_r_c[4]), 
            .I3(GND_net), .O(n11184));
    defparam i9346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13397_bdd_4_lut (.I0(n13397), .I1(\REG.mem_29_3 ), .I2(\REG.mem_28_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11077));
    defparam n13397_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9347_3_lut (.I0(n12842), .I1(n11184), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [14]));
    defparam i9347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9224_3_lut (.I0(n12734), .I1(n13532), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [15]));
    defparam i9224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9636_3_lut (.I0(\REG.mem_48_7 ), .I1(\REG.mem_49_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11474));
    defparam i9636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9637_3_lut (.I0(\REG.mem_50_7 ), .I1(\REG.mem_51_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11475));
    defparam i9637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9667_3_lut (.I0(\REG.mem_54_7 ), .I1(\REG.mem_55_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11505));
    defparam i9667_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i236_237 (.Q(\REG.mem_2_2 ), .C(FIFO_CLK_c), .D(n4947));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9666_3_lut (.I0(\REG.mem_52_7 ), .I1(\REG.mem_53_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11504));
    defparam i9666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10866 (.I0(rd_addr_r_c[2]), .I1(n11068), 
            .I2(n11077), .I3(rd_addr_r_c[3]), .O(n12749));
    defparam rd_addr_r_2__bdd_4_lut_10866.LUT_INIT = 16'he4aa;
    SB_LUT4 i4091_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_34_0 ), .O(n5474));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4091_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12425_bdd_4_lut (.I0(n12425), .I1(\REG.mem_1_13 ), .I2(\REG.mem_0_13 ), 
            .I3(rd_addr_r_c[1]), .O(n11815));
    defparam n12425_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12749_bdd_4_lut (.I0(n12749), .I1(n11065), .I2(n11059), .I3(rd_addr_r_c[3]), 
            .O(n11137));
    defparam n12749_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11375 (.I0(rd_addr_r_c[1]), .I1(n11555), 
            .I2(n11556), .I3(rd_addr_r_c[2]), .O(n13391));
    defparam rd_addr_r_1__bdd_4_lut_11375.LUT_INIT = 16'he4aa;
    SB_LUT4 i9678_3_lut (.I0(\REG.mem_48_10 ), .I1(\REG.mem_49_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11516));
    defparam i9678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9679_3_lut (.I0(\REG.mem_50_10 ), .I1(\REG.mem_51_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11517));
    defparam i9679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10871 (.I0(rd_addr_r_c[1]), .I1(n11870), 
            .I2(n11871), .I3(rd_addr_r_c[2]), .O(n12743));
    defparam rd_addr_r_1__bdd_4_lut_10871.LUT_INIT = 16'he4aa;
    SB_LUT4 n13391_bdd_4_lut (.I0(n13391), .I1(n11541), .I2(n11540), .I3(rd_addr_r_c[2]), 
            .O(n13394));
    defparam n13391_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i6_2_lut_4_lut (.I0(wr_grey_sync_r[6]), 
            .I1(wr_addr_p1_w[6]), .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[5] ), 
            .O(wr_grey_w[5]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i6_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 n12743_bdd_4_lut (.I0(n12743), .I1(n11868), .I2(n11867), .I3(rd_addr_r_c[2]), 
            .O(n12746));
    defparam n12743_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9604_3_lut (.I0(\REG.mem_22_8 ), .I1(\REG.mem_23_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11442));
    defparam i9604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10563 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_9 ), 
            .I2(\REG.mem_59_9 ), .I3(rd_addr_r_c[1]), .O(n12419));
    defparam rd_addr_r_0__bdd_4_lut_10563.LUT_INIT = 16'he4aa;
    SB_LUT4 i9603_3_lut (.I0(\REG.mem_20_8 ), .I1(\REG.mem_21_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11441));
    defparam i9603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11370 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_5 ), 
            .I2(\REG.mem_27_5 ), .I3(rd_addr_r_c[1]), .O(n13385));
    defparam rd_addr_r_0__bdd_4_lut_11370.LUT_INIT = 16'he4aa;
    SB_LUT4 i4289_2_lut_4_lut (.I0(wr_grey_sync_r[6]), .I1(wr_addr_p1_w[6]), 
            .I2(wr_sig_mv_w), .I3(reset_per_frame), .O(n5672));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i4289_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 n13385_bdd_4_lut (.I0(n13385), .I1(\REG.mem_25_5 ), .I2(\REG.mem_24_5 ), 
            .I3(rd_addr_r_c[1]), .O(n13388));
    defparam n13385_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR rd_grey_sync_r__i0 (.Q(\rd_grey_sync_r[0] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[0]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10836 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_15 ), 
            .I2(\REG.mem_27_15 ), .I3(rd_addr_r_c[1]), .O(n12737));
    defparam rd_addr_r_0__bdd_4_lut_10836.LUT_INIT = 16'he4aa;
    SB_LUT4 n12737_bdd_4_lut (.I0(n12737), .I1(\REG.mem_25_15 ), .I2(\REG.mem_24_15 ), 
            .I3(rd_addr_r_c[1]), .O(n12740));
    defparam n12737_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9730_3_lut (.I0(n12326), .I1(n13850), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11568));
    defparam i9730_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i233_234 (.Q(\REG.mem_2_1 ), .C(FIFO_CLK_c), .D(n4946));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9729_3_lut (.I0(n12542), .I1(n12362), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11567));
    defparam i9729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11360 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_12 ), 
            .I2(\REG.mem_15_12 ), .I3(rd_addr_r_c[1]), .O(n13379));
    defparam rd_addr_r_0__bdd_4_lut_11360.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10861 (.I0(rd_addr_r_c[3]), .I1(n12650), 
            .I2(n11016), .I3(rd_addr_r_c[4]), .O(n12731));
    defparam rd_addr_r_3__bdd_4_lut_10861.LUT_INIT = 16'he4aa;
    SB_DFFSS empty_ext_r_124 (.Q(DEBUG_3_c), .C(SLM_CLK_c), .D(empty_nxt_c_N_629), 
            .S(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_LUT4 n13379_bdd_4_lut (.I0(n13379), .I1(\REG.mem_13_12 ), .I2(\REG.mem_12_12 ), 
            .I3(rd_addr_r_c[1]), .O(n13382));
    defparam n13379_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i230_231 (.Q(\REG.mem_2_0 ), .C(FIFO_CLK_c), .D(n4945));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFSR wr_grey_sync_r__i0 (.Q(wr_grey_sync_r[0]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[0]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFF i38_39 (.Q(\REG.mem_0_0 ), .C(FIFO_CLK_c), .D(n4944));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11440 (.I0(rd_addr_r_c[3]), .I1(n13070), 
            .I2(n11586), .I3(rd_addr_r_c[4]), .O(n13373));
    defparam rd_addr_r_3__bdd_4_lut_11440.LUT_INIT = 16'he4aa;
    SB_DFF i41_42 (.Q(\REG.mem_0_1 ), .C(FIFO_CLK_c), .D(n4943));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFS \aempty_flag_impl.ae_flag_ext_r_130  (.Q(dc32_fifo_almost_empty), 
            .C(SLM_CLK_c), .D(\aempty_flag_impl.ae_flag_nxt_w ), .S(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(669[37] 672[40])
    SB_LUT4 i9715_3_lut (.I0(n13154), .I1(n12656), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11553));
    defparam i9715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12731_bdd_4_lut (.I0(n12731), .I1(n11952), .I2(n11951), .I3(rd_addr_r_c[4]), 
            .O(n12734));
    defparam n12731_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13373_bdd_4_lut (.I0(n13373), .I1(n11562), .I2(n13052), .I3(rd_addr_r_c[4]), 
            .O(n13376));
    defparam n13373_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11355 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_1 ), 
            .I2(\REG.mem_7_1 ), .I3(rd_addr_r_c[1]), .O(n13367));
    defparam rd_addr_r_0__bdd_4_lut_11355.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10831 (.I0(rd_addr_r_c[2]), .I1(n11623), 
            .I2(n11632), .I3(rd_addr_r_c[3]), .O(n12725));
    defparam rd_addr_r_2__bdd_4_lut_10831.LUT_INIT = 16'he4aa;
    SB_LUT4 n13367_bdd_4_lut (.I0(n13367), .I1(\REG.mem_5_1 ), .I2(\REG.mem_4_1 ), 
            .I3(rd_addr_r_c[1]), .O(n11230));
    defparam n13367_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12419_bdd_4_lut (.I0(n12419), .I1(\REG.mem_57_9 ), .I2(\REG.mem_56_9 ), 
            .I3(rd_addr_r_c[1]), .O(n12422));
    defparam n12419_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12725_bdd_4_lut (.I0(n12725), .I1(n11611), .I2(n11608), .I3(rd_addr_r_c[3]), 
            .O(n11743));
    defparam n12725_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9181_3_lut (.I0(n13778), .I1(n13754), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11019));
    defparam i9181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10826 (.I0(rd_addr_r_c[1]), .I1(n11894), 
            .I2(n11895), .I3(rd_addr_r_c[2]), .O(n12719));
    defparam rd_addr_r_1__bdd_4_lut_10826.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11345 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_3 ), 
            .I2(\REG.mem_35_3 ), .I3(rd_addr_r_c[1]), .O(n13361));
    defparam rd_addr_r_0__bdd_4_lut_11345.LUT_INIT = 16'he4aa;
    SB_LUT4 n13361_bdd_4_lut (.I0(n13361), .I1(\REG.mem_33_3 ), .I2(\REG.mem_32_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11080));
    defparam n13361_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12719_bdd_4_lut (.I0(n12719), .I1(n11883), .I2(n11882), .I3(rd_addr_r_c[2]), 
            .O(n12722));
    defparam n12719_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11340 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_1 ), 
            .I2(\REG.mem_47_1 ), .I3(rd_addr_r_c[1]), .O(n13355));
    defparam rd_addr_r_0__bdd_4_lut_11340.LUT_INIT = 16'he4aa;
    SB_LUT4 n13355_bdd_4_lut (.I0(n13355), .I1(\REG.mem_45_1 ), .I2(\REG.mem_44_1 ), 
            .I3(rd_addr_r_c[1]), .O(n13358));
    defparam n13355_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10047_3_lut (.I0(\REG.mem_24_2 ), .I1(\REG.mem_25_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11885));
    defparam i10047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10806 (.I0(rd_addr_r_c[1]), .I1(n11864), 
            .I2(n11865), .I3(rd_addr_r_c[2]), .O(n12713));
    defparam rd_addr_r_1__bdd_4_lut_10806.LUT_INIT = 16'he4aa;
    SB_LUT4 i3825_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_17_15 ), .O(n5208));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3825_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3824_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_17_14 ), .O(n5207));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3824_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10048_3_lut (.I0(\REG.mem_26_2 ), .I1(\REG.mem_27_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11886));
    defparam i10048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3823_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_17_13 ), .O(n5206));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3823_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11335 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_11 ), 
            .I2(\REG.mem_3_11 ), .I3(rd_addr_r_c[1]), .O(n13349));
    defparam rd_addr_r_0__bdd_4_lut_11335.LUT_INIT = 16'he4aa;
    SB_DFF i44_45 (.Q(\REG.mem_0_2 ), .C(FIFO_CLK_c), .D(n4941));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13349_bdd_4_lut (.I0(n13349), .I1(\REG.mem_1_11 ), .I2(\REG.mem_0_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11608));
    defparam n13349_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12713_bdd_4_lut (.I0(n12713), .I1(n11856), .I2(n11855), .I3(rd_addr_r_c[2]), 
            .O(n12716));
    defparam n12713_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10060_3_lut (.I0(\REG.mem_30_2 ), .I1(\REG.mem_31_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11898));
    defparam i10060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10059_3_lut (.I0(\REG.mem_28_2 ), .I1(\REG.mem_29_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11897));
    defparam i10059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10821 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_12 ), 
            .I2(\REG.mem_51_12 ), .I3(rd_addr_r_c[1]), .O(n12707));
    defparam rd_addr_r_0__bdd_4_lut_10821.LUT_INIT = 16'he4aa;
    SB_LUT4 i3822_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_17_12 ), .O(n5205));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3822_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11330 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_11 ), 
            .I2(\REG.mem_7_11 ), .I3(rd_addr_r_c[1]), .O(n13343));
    defparam rd_addr_r_0__bdd_4_lut_11330.LUT_INIT = 16'he4aa;
    SB_LUT4 n13343_bdd_4_lut (.I0(n13343), .I1(\REG.mem_5_11 ), .I2(\REG.mem_4_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11611));
    defparam n13343_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3821_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_17_11 ), .O(n5204));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3821_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12305_bdd_4_lut (.I0(n12305), .I1(n11232), .I2(n11231), .I3(rd_addr_r_c[2]), 
            .O(n12308));
    defparam n12305_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12707_bdd_4_lut (.I0(n12707), .I1(\REG.mem_49_12 ), .I2(\REG.mem_48_12 ), 
            .I3(rd_addr_r_c[1]), .O(n12710));
    defparam n12707_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10474 (.I0(rd_addr_r_c[2]), .I1(n11965), 
            .I2(n11971), .I3(rd_addr_r_c[3]), .O(n12311));
    defparam rd_addr_r_2__bdd_4_lut_10474.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10479 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_4 ), 
            .I2(\REG.mem_3_4 ), .I3(rd_addr_r_c[1]), .O(n12299));
    defparam rd_addr_r_0__bdd_4_lut_10479.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10796 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_8 ), 
            .I2(\REG.mem_15_8 ), .I3(rd_addr_r_c[1]), .O(n12701));
    defparam rd_addr_r_0__bdd_4_lut_10796.LUT_INIT = 16'he4aa;
    SB_LUT4 i10020_3_lut (.I0(\REG.mem_8_14 ), .I1(\REG.mem_9_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11858));
    defparam i10020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3820_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_17_10 ), .O(n5203));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3820_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10021_3_lut (.I0(\REG.mem_10_14 ), .I1(\REG.mem_11_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11859));
    defparam i10021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11325 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_6 ), 
            .I2(\REG.mem_63_6 ), .I3(rd_addr_r_c[1]), .O(n13337));
    defparam rd_addr_r_0__bdd_4_lut_11325.LUT_INIT = 16'he4aa;
    SB_DFF i47_48 (.Q(\REG.mem_0_3 ), .C(FIFO_CLK_c), .D(n4940));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12701_bdd_4_lut (.I0(n12701), .I1(\REG.mem_13_8 ), .I2(\REG.mem_12_8 ), 
            .I3(rd_addr_r_c[1]), .O(n12704));
    defparam n12701_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10024_3_lut (.I0(\REG.mem_14_14 ), .I1(\REG.mem_15_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11862));
    defparam i10024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10816 (.I0(rd_addr_r_c[3]), .I1(n11012), 
            .I2(n12470), .I3(rd_addr_r_c[4]), .O(n12695));
    defparam rd_addr_r_3__bdd_4_lut_10816.LUT_INIT = 16'he4aa;
    SB_LUT4 i3819_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_17_9 ), .O(n5202));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3819_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3818_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_17_8 ), .O(n5201));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3818_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10558 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_1 ), 
            .I2(\REG.mem_3_1 ), .I3(rd_addr_r_c[1]), .O(n12413));
    defparam rd_addr_r_0__bdd_4_lut_10558.LUT_INIT = 16'he4aa;
    SB_LUT4 i3817_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_17_7 ), .O(n5200));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3817_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12695_bdd_4_lut (.I0(n12695), .I1(n11010), .I2(n11009), .I3(rd_addr_r_c[4]), 
            .O(n12698));
    defparam n12695_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10023_3_lut (.I0(\REG.mem_12_14 ), .I1(\REG.mem_13_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11861));
    defparam i10023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10801 (.I0(rd_addr_r_c[1]), .I1(n11852), 
            .I2(n11853), .I3(rd_addr_r_c[2]), .O(n12689));
    defparam rd_addr_r_1__bdd_4_lut_10801.LUT_INIT = 16'he4aa;
    SB_LUT4 n13337_bdd_4_lut (.I0(n13337), .I1(\REG.mem_61_6 ), .I2(\REG.mem_60_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11614));
    defparam n13337_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3816_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_17_6 ), .O(n5199));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3816_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12689_bdd_4_lut (.I0(n12689), .I1(n11850), .I2(n11849), .I3(rd_addr_r_c[2]), 
            .O(n12692));
    defparam n12689_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3815_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_17_5 ), .O(n5198));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3815_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3814_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_17_4 ), .O(n5197));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3814_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11350 (.I0(rd_addr_r_c[3]), .I1(n13076), 
            .I2(n11595), .I3(rd_addr_r_c[4]), .O(n13331));
    defparam rd_addr_r_3__bdd_4_lut_11350.LUT_INIT = 16'he4aa;
    SB_LUT4 n13331_bdd_4_lut (.I0(n13331), .I1(n11583), .I2(n13064), .I3(rd_addr_r_c[4]), 
            .O(n13334));
    defparam n13331_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3813_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_17_3 ), .O(n5196));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3813_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10791 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_8 ), 
            .I2(\REG.mem_43_8 ), .I3(rd_addr_r_c[1]), .O(n12683));
    defparam rd_addr_r_0__bdd_4_lut_10791.LUT_INIT = 16'he4aa;
    SB_LUT4 i3812_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_17_2 ), .O(n5195));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3812_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3811_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_17_1 ), .O(n5194));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3811_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11365 (.I0(rd_addr_r_c[1]), .I1(n11171), 
            .I2(n11172), .I3(rd_addr_r_c[2]), .O(n13325));
    defparam rd_addr_r_1__bdd_4_lut_11365.LUT_INIT = 16'he4aa;
    SB_LUT4 n13325_bdd_4_lut (.I0(n13325), .I1(n11169), .I2(n11168), .I3(rd_addr_r_c[2]), 
            .O(n11250));
    defparam n13325_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12683_bdd_4_lut (.I0(n12683), .I1(\REG.mem_41_8 ), .I2(\REG.mem_40_8 ), 
            .I3(rd_addr_r_c[1]), .O(n12686));
    defparam n12683_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3810_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_17_0 ), .O(n5193));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3810_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_addr_r_6__I_0_135_i6_3_lut (.I0(wr_addr_r[5]), .I1(wr_addr_p1_w[5]), 
            .I2(wr_sig_mv_w), .I3(GND_net), .O(\wr_addr_nxt_c[5] ));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_6__I_0_135_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10782 (.I0(rd_addr_r_c[1]), .I1(n11948), 
            .I2(n11949), .I3(rd_addr_r_c[2]), .O(n12677));
    defparam rd_addr_r_1__bdd_4_lut_10782.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11320 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_12 ), 
            .I2(\REG.mem_19_12 ), .I3(rd_addr_r_c[1]), .O(n13319));
    defparam rd_addr_r_0__bdd_4_lut_11320.LUT_INIT = 16'he4aa;
    SB_LUT4 n12413_bdd_4_lut (.I0(n12413), .I1(\REG.mem_1_1 ), .I2(\REG.mem_0_1 ), 
            .I3(rd_addr_r_c[1]), .O(n12416));
    defparam n12413_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3857_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_19_15 ), .O(n5240));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3857_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13319_bdd_4_lut (.I0(n13319), .I1(\REG.mem_17_12 ), .I2(\REG.mem_16_12 ), 
            .I3(rd_addr_r_c[1]), .O(n13322));
    defparam n13319_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3856_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_19_14 ), .O(n5239));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3856_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3855_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_19_13 ), .O(n5238));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3855_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12677_bdd_4_lut (.I0(n12677), .I1(n11943), .I2(n11942), .I3(rd_addr_r_c[2]), 
            .O(n12680));
    defparam n12677_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3854_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_19_12 ), .O(n5237));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3854_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3853_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_19_11 ), .O(n5236));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3853_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3852_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_19_10 ), .O(n5235));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3852_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3851_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_19_9 ), .O(n5234));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3851_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3850_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_19_8 ), .O(n5233));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3850_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10772 (.I0(rd_addr_r_c[1]), .I1(n11909), 
            .I2(n11910), .I3(rd_addr_r_c[2]), .O(n12671));
    defparam rd_addr_r_1__bdd_4_lut_10772.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11310 (.I0(rd_addr_r_c[1]), .I1(n11198), 
            .I2(n11199), .I3(rd_addr_r_c[2]), .O(n13313));
    defparam rd_addr_r_1__bdd_4_lut_11310.LUT_INIT = 16'he4aa;
    SB_LUT4 i3849_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_19_7 ), .O(n5232));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3849_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12671_bdd_4_lut (.I0(n12671), .I1(n11907), .I2(n11906), .I3(rd_addr_r_c[2]), 
            .O(n12674));
    defparam n12671_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3848_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_19_6 ), .O(n5231));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3848_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10777 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_15 ), 
            .I2(\REG.mem_31_15 ), .I3(rd_addr_r_c[1]), .O(n12665));
    defparam rd_addr_r_0__bdd_4_lut_10777.LUT_INIT = 16'he4aa;
    SB_LUT4 n13313_bdd_4_lut (.I0(n13313), .I1(n11193), .I2(n11192), .I3(rd_addr_r_c[2]), 
            .O(n11256));
    defparam n13313_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3847_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_19_5 ), .O(n5230));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3847_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3846_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_19_4 ), .O(n5229));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3846_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3845_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_19_3 ), .O(n5228));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3845_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12665_bdd_4_lut (.I0(n12665), .I1(\REG.mem_29_15 ), .I2(\REG.mem_28_15 ), 
            .I3(rd_addr_r_c[1]), .O(n12668));
    defparam n12665_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11305 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_3 ), 
            .I2(\REG.mem_39_3 ), .I3(rd_addr_r_c[1]), .O(n13307));
    defparam rd_addr_r_0__bdd_4_lut_11305.LUT_INIT = 16'he4aa;
    SB_LUT4 n13307_bdd_4_lut (.I0(n13307), .I1(\REG.mem_37_3 ), .I2(\REG.mem_36_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11086));
    defparam n13307_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10811 (.I0(rd_addr_r_c[2]), .I1(n11656), 
            .I2(n11668), .I3(rd_addr_r_c[3]), .O(n12659));
    defparam rd_addr_r_2__bdd_4_lut_10811.LUT_INIT = 16'he4aa;
    SB_LUT4 n12659_bdd_4_lut (.I0(n12659), .I1(n11653), .I2(n11644), .I3(rd_addr_r_c[3]), 
            .O(n11755));
    defparam n12659_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3844_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_19_2 ), .O(n5227));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3844_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11295 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_3 ), 
            .I2(\REG.mem_43_3 ), .I3(rd_addr_r_c[1]), .O(n13301));
    defparam rd_addr_r_0__bdd_4_lut_11295.LUT_INIT = 16'he4aa;
    SB_LUT4 i3843_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_19_1 ), .O(n5226));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3843_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10762 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_7 ), 
            .I2(\REG.mem_15_7 ), .I3(rd_addr_r_c[1]), .O(n12653));
    defparam rd_addr_r_0__bdd_4_lut_10762.LUT_INIT = 16'he4aa;
    SB_LUT4 n12653_bdd_4_lut (.I0(n12653), .I1(\REG.mem_13_7 ), .I2(\REG.mem_12_7 ), 
            .I3(rd_addr_r_c[1]), .O(n12656));
    defparam n12653_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13301_bdd_4_lut (.I0(n13301), .I1(\REG.mem_41_3 ), .I2(\REG.mem_40_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11089));
    defparam n13301_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10767 (.I0(rd_addr_r_c[1]), .I1(n11714), 
            .I2(n11715), .I3(rd_addr_r_c[2]), .O(n12647));
    defparam rd_addr_r_1__bdd_4_lut_10767.LUT_INIT = 16'he4aa;
    SB_LUT4 i3842_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_19_0 ), .O(n5225));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3842_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12647_bdd_4_lut (.I0(n12647), .I1(n11694), .I2(n11693), .I3(rd_addr_r_c[2]), 
            .O(n12650));
    defparam n12647_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11290 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_0 ), 
            .I2(\REG.mem_59_0 ), .I3(rd_addr_r_c[1]), .O(n13295));
    defparam rd_addr_r_0__bdd_4_lut_11290.LUT_INIT = 16'he4aa;
    SB_LUT4 n13295_bdd_4_lut (.I0(n13295), .I1(\REG.mem_57_0 ), .I2(\REG.mem_56_0 ), 
            .I3(rd_addr_r_c[1]), .O(n13298));
    defparam n13295_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10747 (.I0(rd_addr_r_c[1]), .I1(n11681), 
            .I2(n11682), .I3(rd_addr_r_c[2]), .O(n12641));
    defparam rd_addr_r_1__bdd_4_lut_10747.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11285 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_11 ), 
            .I2(\REG.mem_11_11 ), .I3(rd_addr_r_c[1]), .O(n13289));
    defparam rd_addr_r_0__bdd_4_lut_11285.LUT_INIT = 16'he4aa;
    SB_LUT4 n12641_bdd_4_lut (.I0(n12641), .I1(n11637), .I2(n11636), .I3(rd_addr_r_c[2]), 
            .O(n12644));
    defparam n12641_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13289_bdd_4_lut (.I0(n13289), .I1(\REG.mem_9_11 ), .I2(\REG.mem_8_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11623));
    defparam n13289_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10553 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_12 ), 
            .I2(\REG.mem_63_12 ), .I3(rd_addr_r_c[1]), .O(n12407));
    defparam rd_addr_r_0__bdd_4_lut_10553.LUT_INIT = 16'he4aa;
    SB_LUT4 i3873_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_20_15 ), .O(n5256));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3873_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3872_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_20_14 ), .O(n5255));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3872_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3871_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_20_13 ), .O(n5254));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3871_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3870_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_20_12 ), .O(n5253));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3870_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3869_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_20_11 ), .O(n5252));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3869_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3868_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_20_10 ), .O(n5251));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3868_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10757 (.I0(rd_addr_r_c[2]), .I1(n10993), 
            .I2(n10996), .I3(rd_addr_r_c[3]), .O(n12635));
    defparam rd_addr_r_2__bdd_4_lut_10757.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11315 (.I0(rd_addr_r_c[3]), .I1(n12716), 
            .I2(n11049), .I3(rd_addr_r_c[4]), .O(n13283));
    defparam rd_addr_r_3__bdd_4_lut_11315.LUT_INIT = 16'he4aa;
    SB_LUT4 n12635_bdd_4_lut (.I0(n12635), .I1(n12016), .I2(n12010), .I3(rd_addr_r_c[3]), 
            .O(n12638));
    defparam n12635_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3867_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_20_9 ), .O(n5250));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3867_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10752 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_12 ), 
            .I2(\REG.mem_55_12 ), .I3(rd_addr_r_c[1]), .O(n12629));
    defparam rd_addr_r_0__bdd_4_lut_10752.LUT_INIT = 16'he4aa;
    SB_LUT4 n13283_bdd_4_lut (.I0(n13283), .I1(n11004), .I2(n12644), .I3(rd_addr_r_c[4]), 
            .O(n13286));
    defparam n13283_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12629_bdd_4_lut (.I0(n12629), .I1(\REG.mem_53_12 ), .I2(\REG.mem_52_12 ), 
            .I3(rd_addr_r_c[1]), .O(n12632));
    defparam n12629_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11300 (.I0(rd_addr_r_c[1]), .I1(n11219), 
            .I2(n11220), .I3(rd_addr_r_c[2]), .O(n13277));
    defparam rd_addr_r_1__bdd_4_lut_11300.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10732 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_15 ), 
            .I2(\REG.mem_35_15 ), .I3(rd_addr_r_c[1]), .O(n12623));
    defparam rd_addr_r_0__bdd_4_lut_10732.LUT_INIT = 16'he4aa;
    SB_LUT4 n12623_bdd_4_lut (.I0(n12623), .I1(\REG.mem_33_15 ), .I2(\REG.mem_32_15 ), 
            .I3(rd_addr_r_c[1]), .O(n12626));
    defparam n12623_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13277_bdd_4_lut (.I0(n13277), .I1(n11217), .I2(n11216), .I3(rd_addr_r_c[2]), 
            .O(n11259));
    defparam n13277_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11280 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_15 ), 
            .I2(\REG.mem_3_15 ), .I3(rd_addr_r_c[1]), .O(n13271));
    defparam rd_addr_r_0__bdd_4_lut_11280.LUT_INIT = 16'he4aa;
    SB_LUT4 i3866_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_20_8 ), .O(n5249));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3866_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3865_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_20_7 ), .O(n5248));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3865_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_addr_r_6__I_0_135_i4_3_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_w[3]), 
            .I2(wr_sig_mv_w), .I3(GND_net), .O(\wr_addr_nxt_c[3] ));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_6__I_0_135_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13271_bdd_4_lut (.I0(n13271), .I1(\REG.mem_1_15 ), .I2(\REG.mem_0_15 ), 
            .I3(rd_addr_r_c[1]), .O(n13274));
    defparam n13271_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i50_51 (.Q(\REG.mem_0_4 ), .C(FIFO_CLK_c), .D(n4935));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10727 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_9 ), 
            .I2(\REG.mem_51_9 ), .I3(rd_addr_r_c[1]), .O(n12617));
    defparam rd_addr_r_0__bdd_4_lut_10727.LUT_INIT = 16'he4aa;
    SB_DFF i53_54 (.Q(\REG.mem_0_5 ), .C(FIFO_CLK_c), .D(n4934));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12617_bdd_4_lut (.I0(n12617), .I1(\REG.mem_49_9 ), .I2(\REG.mem_48_9 ), 
            .I3(rd_addr_r_c[1]), .O(n12620));
    defparam n12617_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3864_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_20_6 ), .O(n5247));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3864_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3863_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_20_5 ), .O(n5246));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3863_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12299_bdd_4_lut (.I0(n12299), .I1(\REG.mem_1_4 ), .I2(\REG.mem_0_4 ), 
            .I3(rd_addr_r_c[1]), .O(n12302));
    defparam n12299_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10460 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_8 ), 
            .I2(\REG.mem_47_8 ), .I3(rd_addr_r_c[1]), .O(n12293));
    defparam rd_addr_r_0__bdd_4_lut_10460.LUT_INIT = 16'he4aa;
    SB_LUT4 i3862_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_20_4 ), .O(n5245));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3862_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3861_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_20_3 ), .O(n5244));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3861_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11265 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_3 ), 
            .I2(\REG.mem_47_3 ), .I3(rd_addr_r_c[1]), .O(n13265));
    defparam rd_addr_r_0__bdd_4_lut_11265.LUT_INIT = 16'he4aa;
    SB_LUT4 n12293_bdd_4_lut (.I0(n12293), .I1(\REG.mem_45_8 ), .I2(\REG.mem_44_8 ), 
            .I3(rd_addr_r_c[1]), .O(n12296));
    defparam n12293_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12335_bdd_4_lut (.I0(n12335), .I1(\REG.mem_17_2 ), .I2(\REG.mem_16_2 ), 
            .I3(rd_addr_r_c[1]), .O(n12338));
    defparam n12335_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10489 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_9 ), 
            .I2(\REG.mem_11_9 ), .I3(rd_addr_r_c[1]), .O(n12329));
    defparam rd_addr_r_0__bdd_4_lut_10489.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10737 (.I0(rd_addr_r_c[2]), .I1(n11692), 
            .I2(n11701), .I3(rd_addr_r_c[3]), .O(n12611));
    defparam rd_addr_r_2__bdd_4_lut_10737.LUT_INIT = 16'he4aa;
    SB_LUT4 n13265_bdd_4_lut (.I0(n13265), .I1(\REG.mem_45_3 ), .I2(\REG.mem_44_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11104));
    defparam n13265_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3860_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_20_2 ), .O(n5243));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3860_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3859_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_20_1 ), .O(n5242));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3859_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12323_bdd_4_lut (.I0(n12323), .I1(\REG.mem_25_7 ), .I2(\REG.mem_24_7 ), 
            .I3(rd_addr_r_c[1]), .O(n12326));
    defparam n12323_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11260 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_12 ), 
            .I2(\REG.mem_23_12 ), .I3(rd_addr_r_c[1]), .O(n13259));
    defparam rd_addr_r_0__bdd_4_lut_11260.LUT_INIT = 16'he4aa;
    SB_LUT4 i3858_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_20_0 ), .O(n5241));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3858_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12611_bdd_4_lut (.I0(n12611), .I1(n11677), .I2(n11674), .I3(rd_addr_r_c[3]), 
            .O(n11764));
    defparam n12611_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10587 (.I0(rd_addr_r_c[2]), .I1(n11158), 
            .I2(n11176), .I3(rd_addr_r_c[3]), .O(n12317));
    defparam rd_addr_r_2__bdd_4_lut_10587.LUT_INIT = 16'he4aa;
    SB_LUT4 i3890_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_21_15 ), .O(n5273));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3890_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13259_bdd_4_lut (.I0(n13259), .I1(\REG.mem_21_12 ), .I2(\REG.mem_20_12 ), 
            .I3(rd_addr_r_c[1]), .O(n13262));
    defparam n13259_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12407_bdd_4_lut (.I0(n12407), .I1(\REG.mem_61_12 ), .I2(\REG.mem_60_12 ), 
            .I3(rd_addr_r_c[1]), .O(n12410));
    defparam n12407_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12311_bdd_4_lut (.I0(n12311), .I1(n11959), .I2(n11815), .I3(rd_addr_r_c[3]), 
            .O(n12314));
    defparam n12311_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3889_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_21_14 ), .O(n5272));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3889_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3888_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_21_13 ), .O(n5271));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3888_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10494 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_2 ), 
            .I2(\REG.mem_19_2 ), .I3(rd_addr_r_c[1]), .O(n12335));
    defparam rd_addr_r_0__bdd_4_lut_10494.LUT_INIT = 16'he4aa;
    SB_LUT4 i3887_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_21_12 ), .O(n5270));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3887_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3886_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_21_11 ), .O(n5269));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3886_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i5_1_lut (.I0(rd_addr_r_c[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3885_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_21_10 ), .O(n5268));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3885_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3884_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_21_9 ), .O(n5267));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3884_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10722 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_0 ), 
            .I2(\REG.mem_39_0 ), .I3(rd_addr_r_c[1]), .O(n12605));
    defparam rd_addr_r_0__bdd_4_lut_10722.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10469 (.I0(rd_addr_r_c[2]), .I1(n11455), 
            .I2(n11488), .I3(rd_addr_r_c[3]), .O(n12287));
    defparam rd_addr_r_2__bdd_4_lut_10469.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11255 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_13 ), 
            .I2(\REG.mem_31_13 ), .I3(rd_addr_r_c[1]), .O(n13253));
    defparam rd_addr_r_0__bdd_4_lut_11255.LUT_INIT = 16'he4aa;
    SB_LUT4 n12605_bdd_4_lut (.I0(n12605), .I1(\REG.mem_37_0 ), .I2(\REG.mem_36_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11332));
    defparam n12605_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13253_bdd_4_lut (.I0(n13253), .I1(\REG.mem_29_13 ), .I2(\REG.mem_28_13 ), 
            .I3(rd_addr_r_c[1]), .O(n13256));
    defparam n13253_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3883_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_21_8 ), .O(n5266));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3883_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10717 (.I0(rd_addr_r_c[2]), .I1(n11722), 
            .I2(n11737), .I3(rd_addr_r_c[3]), .O(n12599));
    defparam rd_addr_r_2__bdd_4_lut_10717.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11250 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_6 ), 
            .I2(\REG.mem_19_6 ), .I3(rd_addr_r_c[1]), .O(n13247));
    defparam rd_addr_r_0__bdd_4_lut_11250.LUT_INIT = 16'he4aa;
    SB_LUT4 n13247_bdd_4_lut (.I0(n13247), .I1(\REG.mem_17_6 ), .I2(\REG.mem_16_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11110));
    defparam n13247_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3882_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_21_7 ), .O(n5265));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3882_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3881_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_21_6 ), .O(n5264));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3881_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3880_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_21_5 ), .O(n5263));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3880_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3879_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_21_4 ), .O(n5262));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3879_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3878_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_21_3 ), .O(n5261));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3878_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12329_bdd_4_lut (.I0(n12329), .I1(\REG.mem_9_9 ), .I2(\REG.mem_8_9 ), 
            .I3(rd_addr_r_c[1]), .O(n11158));
    defparam n12329_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11245 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_3 ), 
            .I2(\REG.mem_51_3 ), .I3(rd_addr_r_c[1]), .O(n13241));
    defparam rd_addr_r_0__bdd_4_lut_11245.LUT_INIT = 16'he4aa;
    SB_LUT4 n12599_bdd_4_lut (.I0(n12599), .I1(n11719), .I2(n11710), .I3(rd_addr_r_c[3]), 
            .O(n11767));
    defparam n12599_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13241_bdd_4_lut (.I0(n13241), .I1(\REG.mem_49_3 ), .I2(\REG.mem_48_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11113));
    defparam n13241_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3877_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_21_2 ), .O(n5260));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3877_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3876_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_21_1 ), .O(n5259));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3876_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10712 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_0 ), 
            .I2(\REG.mem_43_0 ), .I3(rd_addr_r_c[1]), .O(n12593));
    defparam rd_addr_r_0__bdd_4_lut_10712.LUT_INIT = 16'he4aa;
    SB_LUT4 i3874_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_21_0 ), .O(n5257));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3874_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3906_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_22_15 ), .O(n5289));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3906_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3905_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_22_14 ), .O(n5288));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3905_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3904_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_22_13 ), .O(n5287));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3904_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11270 (.I0(rd_addr_r_c[1]), .I1(n11996), 
            .I2(n11997), .I3(rd_addr_r_c[2]), .O(n13235));
    defparam rd_addr_r_1__bdd_4_lut_11270.LUT_INIT = 16'he4aa;
    SB_LUT4 n12593_bdd_4_lut (.I0(n12593), .I1(\REG.mem_41_0 ), .I2(\REG.mem_40_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11335));
    defparam n12593_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13235_bdd_4_lut (.I0(n13235), .I1(n11991), .I2(n11990), .I3(rd_addr_r_c[2]), 
            .O(n13238));
    defparam n13235_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3903_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_22_12 ), .O(n5286));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3903_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3902_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_22_11 ), .O(n5285));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3902_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3901_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_22_10 ), .O(n5284));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3901_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3900_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_22_9 ), .O(n5283));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3900_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3899_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_22_8 ), .O(n5282));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3899_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3898_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_22_7 ), .O(n5281));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3898_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3897_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_22_6 ), .O(n5280));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3897_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3896_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_22_5 ), .O(n5279));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3896_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3895_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_22_4 ), .O(n5278));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3895_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3894_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_22_3 ), .O(n5277));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3894_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3893_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_22_2 ), .O(n5276));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3893_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11240 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_11 ), 
            .I2(\REG.mem_15_11 ), .I3(rd_addr_r_c[1]), .O(n13229));
    defparam rd_addr_r_0__bdd_4_lut_11240.LUT_INIT = 16'he4aa;
    SB_LUT4 i3892_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_22_1 ), .O(n5275));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3892_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13229_bdd_4_lut (.I0(n13229), .I1(\REG.mem_13_11 ), .I2(\REG.mem_12_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11632));
    defparam n13229_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3891_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_22_0 ), .O(n5274));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3891_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3946_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_24_15 ), .O(n5329));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3946_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_10622 (.I0(rd_addr_r_c[4]), .I1(n11728), 
            .I2(n11785), .I3(rd_addr_r_c[5]), .O(n12401));
    defparam rd_addr_r_4__bdd_4_lut_10622.LUT_INIT = 16'he4aa;
    SB_LUT4 i3945_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_24_14 ), .O(n5328));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3945_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3944_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_24_13 ), .O(n5327));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3944_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12401_bdd_4_lut (.I0(n12401), .I1(n11704), .I2(n11659), .I3(rd_addr_r_c[5]), 
            .O(\REG.out_raw_31__N_559 [6]));
    defparam n12401_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3943_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_24_12 ), .O(n5326));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3943_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11230 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_13 ), 
            .I2(\REG.mem_59_13 ), .I3(rd_addr_r_c[1]), .O(n13223));
    defparam rd_addr_r_0__bdd_4_lut_11230.LUT_INIT = 16'he4aa;
    SB_LUT4 i3942_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_24_11 ), .O(n5325));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3942_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10702 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_5 ), 
            .I2(\REG.mem_39_5 ), .I3(rd_addr_r_c[1]), .O(n12581));
    defparam rd_addr_r_0__bdd_4_lut_10702.LUT_INIT = 16'he4aa;
    SB_LUT4 n12581_bdd_4_lut (.I0(n12581), .I1(\REG.mem_37_5 ), .I2(\REG.mem_36_5 ), 
            .I3(rd_addr_r_c[1]), .O(n12584));
    defparam n12581_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13223_bdd_4_lut (.I0(n13223), .I1(\REG.mem_57_13 ), .I2(\REG.mem_56_13 ), 
            .I3(rd_addr_r_c[1]), .O(n13226));
    defparam n13223_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11235 (.I0(rd_addr_r_c[1]), .I1(n11240), 
            .I2(n11241), .I3(rd_addr_r_c[2]), .O(n13217));
    defparam rd_addr_r_1__bdd_4_lut_11235.LUT_INIT = 16'he4aa;
    SB_LUT4 i3941_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_24_10 ), .O(n5324));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3941_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i56_57 (.Q(\REG.mem_0_6 ), .C(FIFO_CLK_c), .D(n4933));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3940_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_24_9 ), .O(n5323));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3940_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \REG.out_buffer__i2  (.Q(\fifo_data_out[2] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n6121));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 n13217_bdd_4_lut (.I0(n13217), .I1(n11238), .I2(n11237), .I3(rd_addr_r_c[2]), 
            .O(n11262));
    defparam n13217_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \REG.out_buffer__i1  (.Q(\fifo_data_out[1] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n6118));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 i3939_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_24_8 ), .O(n5322));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3939_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3938_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_24_7 ), .O(n5321));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3938_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11225 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_1 ), 
            .I2(\REG.mem_51_1 ), .I3(rd_addr_r_c[1]), .O(n13211));
    defparam rd_addr_r_0__bdd_4_lut_11225.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10692 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_9 ), 
            .I2(\REG.mem_7_9 ), .I3(rd_addr_r_c[1]), .O(n12575));
    defparam rd_addr_r_0__bdd_4_lut_10692.LUT_INIT = 16'he4aa;
    SB_LUT4 i3937_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_24_6 ), .O(n5320));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3937_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13211_bdd_4_lut (.I0(n13211), .I1(\REG.mem_49_1 ), .I2(\REG.mem_48_1 ), 
            .I3(rd_addr_r_c[1]), .O(n13214));
    defparam n13211_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF \REG.out_buffer__i3  (.Q(\fifo_data_out[3] ), .C(SLM_CLK_c), 
           .D(n10556));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i4  (.Q(\fifo_data_out[4] ), .C(SLM_CLK_c), 
           .D(n10562));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i4_1_lut (.I0(rd_addr_r_c[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11215 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_11 ), 
            .I2(\REG.mem_19_11 ), .I3(rd_addr_r_c[1]), .O(n13205));
    defparam rd_addr_r_0__bdd_4_lut_11215.LUT_INIT = 16'he4aa;
    SB_LUT4 i4369_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_49_15 ), .O(n5752));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4369_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13205_bdd_4_lut (.I0(n13205), .I1(\REG.mem_17_11 ), .I2(\REG.mem_16_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11644));
    defparam n13205_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9545_3_lut (.I0(n12956), .I1(n12308), .I2(rd_addr_r_c[3]), 
            .I3(GND_net), .O(n11383));
    defparam i9545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4368_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_49_14 ), .O(n5751));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4368_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3936_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_24_5 ), .O(n5319));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3936_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3935_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_24_4 ), .O(n5318));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3935_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3934_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_24_3 ), .O(n5317));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3934_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3933_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_24_2 ), .O(n5316));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3933_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12575_bdd_4_lut (.I0(n12575), .I1(\REG.mem_5_9 ), .I2(\REG.mem_4_9 ), 
            .I3(rd_addr_r_c[1]), .O(n11143));
    defparam n12575_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3932_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_24_1 ), .O(n5315));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3932_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF \REG.out_buffer__i5  (.Q(\fifo_data_out[5] ), .C(SLM_CLK_c), 
           .D(n10564));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 i3924_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_24_0 ), .O(n5307));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3924_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF \REG.out_buffer__i6  (.Q(\fifo_data_out[6] ), .C(SLM_CLK_c), 
           .D(n10566));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i7  (.Q(\fifo_data_out[7] ), .C(SLM_CLK_c), 
           .D(n10568));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i8  (.Q(\fifo_data_out[8] ), .C(SLM_CLK_c), 
           .D(n10570));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i9  (.Q(\fifo_data_out[9] ), .C(SLM_CLK_c), 
           .D(n10572));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i10  (.Q(\fifo_data_out[10] ), .C(SLM_CLK_c), 
           .D(n10574));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i11  (.Q(\fifo_data_out[11] ), .C(SLM_CLK_c), 
           .D(n10576));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 i4367_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_49_13 ), .O(n5750));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4367_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3978_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_26_15 ), .O(n5361));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3978_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4366_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_49_12 ), .O(n5749));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4366_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3977_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_26_14 ), .O(n5360));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3977_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4365_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_49_11 ), .O(n5748));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4365_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11210 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_5 ), 
            .I2(\REG.mem_31_5 ), .I3(rd_addr_r_c[1]), .O(n13199));
    defparam rd_addr_r_0__bdd_4_lut_11210.LUT_INIT = 16'he4aa;
    SB_LUT4 i4364_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_49_10 ), .O(n5747));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4364_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13199_bdd_4_lut (.I0(n13199), .I1(\REG.mem_29_5 ), .I2(\REG.mem_28_5 ), 
            .I3(rd_addr_r_c[1]), .O(n13202));
    defparam n13199_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \REG.out_buffer__i0  (.Q(\fifo_data_out[0] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n6085));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 i4363_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_49_9 ), .O(n5746));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4363_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4362_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_49_8 ), .O(n5745));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4362_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11205 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_12 ), 
            .I2(\REG.mem_27_12 ), .I3(rd_addr_r_c[1]), .O(n13193));
    defparam rd_addr_r_0__bdd_4_lut_11205.LUT_INIT = 16'he4aa;
    SB_LUT4 i3976_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_26_13 ), .O(n5359));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3976_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3975_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_26_12 ), .O(n5358));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3975_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4361_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_49_7 ), .O(n5744));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4361_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13193_bdd_4_lut (.I0(n13193), .I1(\REG.mem_25_12 ), .I2(\REG.mem_24_12 ), 
            .I3(rd_addr_r_c[1]), .O(n13196));
    defparam n13193_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i6_1_lut (.I0(rd_addr_r_c[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10548 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_13 ), 
            .I2(\REG.mem_39_13 ), .I3(rd_addr_r_c[1]), .O(n12395));
    defparam rd_addr_r_0__bdd_4_lut_10548.LUT_INIT = 16'he4aa;
    SB_LUT4 i4360_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_49_6 ), .O(n5743));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4360_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4359_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_49_5 ), .O(n5742));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4359_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3974_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_26_11 ), .O(n5357));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3974_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4358_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_49_4 ), .O(n5741));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4358_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF \REG.out_buffer__i12  (.Q(\fifo_data_out[12] ), .C(SLM_CLK_c), 
           .D(n10578));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i13  (.Q(\fifo_data_out[13] ), .C(SLM_CLK_c), 
           .D(n10580));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF i59_60 (.Q(\REG.mem_0_7 ), .C(FIFO_CLK_c), .D(n4932));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4357_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_49_3 ), .O(n5740));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4357_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wp_sync2_r_6__I_0_143_i1_2_lut (.I0(wp_sync2_r[5]), .I1(wp_sync2_r[6]), 
            .I2(GND_net), .I3(GND_net), .O(wp_sync_w[5]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam wp_sync2_r_6__I_0_143_i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3973_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_26_10 ), .O(n5356));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3973_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3972_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_26_9 ), .O(n5355));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3972_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i7_1_lut (.I0(\rd_addr_r[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3971_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_26_8 ), .O(n5354));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3971_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3970_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_26_7 ), .O(n5353));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3970_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4356_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_49_2 ), .O(n5739));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4356_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3969_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_26_6 ), .O(n5352));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3969_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11200 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_15 ), 
            .I2(\REG.mem_7_15 ), .I3(rd_addr_r_c[1]), .O(n13187));
    defparam rd_addr_r_0__bdd_4_lut_11200.LUT_INIT = 16'he4aa;
    SB_LUT4 i4355_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_49_1 ), .O(n5738));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4355_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3968_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_26_5 ), .O(n5351));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3968_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF wr_addr_r__i1 (.Q(wr_addr_r[1]), .C(FIFO_CLK_c), .D(n6045));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i2 (.Q(wr_addr_r[2]), .C(FIFO_CLK_c), .D(n6044));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i3 (.Q(wr_addr_r[3]), .C(FIFO_CLK_c), .D(n6043));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i4 (.Q(wr_addr_r[4]), .C(FIFO_CLK_c), .D(n6042));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 n13187_bdd_4_lut (.I0(n13187), .I1(\REG.mem_5_15 ), .I2(\REG.mem_4_15 ), 
            .I3(rd_addr_r_c[1]), .O(n13190));
    defparam n13187_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4354_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_49_0 ), .O(n5737));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4354_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11195 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_13 ), 
            .I2(\REG.mem_35_13 ), .I3(rd_addr_r_c[1]), .O(n13181));
    defparam rd_addr_r_0__bdd_4_lut_11195.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10707 (.I0(rd_addr_r_c[2]), .I1(n11335), 
            .I2(n11947), .I3(rd_addr_r_c[3]), .O(n12551));
    defparam rd_addr_r_2__bdd_4_lut_10707.LUT_INIT = 16'he4aa;
    SB_DFF wr_addr_r__i5 (.Q(wr_addr_r[5]), .C(FIFO_CLK_c), .D(n6024));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF i6131_6132 (.Q(\REG.mem_63_15 ), .C(FIFO_CLK_c), .D(n6021));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6128_6129 (.Q(\REG.mem_63_14 ), .C(FIFO_CLK_c), .D(n6020));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6125_6126 (.Q(\REG.mem_63_13 ), .C(FIFO_CLK_c), .D(n6019));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6122_6123 (.Q(\REG.mem_63_12 ), .C(FIFO_CLK_c), .D(n6018));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i62_63 (.Q(\REG.mem_0_8 ), .C(FIFO_CLK_c), .D(n4931));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12551_bdd_4_lut (.I0(n12551), .I1(n11332), .I2(n11320), .I3(rd_addr_r_c[3]), 
            .O(n12554));
    defparam n12551_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13181_bdd_4_lut (.I0(n13181), .I1(\REG.mem_33_13 ), .I2(\REG.mem_32_13 ), 
            .I3(rd_addr_r_c[1]), .O(n13184));
    defparam n13181_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11190 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_6 ), 
            .I2(\REG.mem_27_6 ), .I3(rd_addr_r_c[1]), .O(n13175));
    defparam rd_addr_r_0__bdd_4_lut_11190.LUT_INIT = 16'he4aa;
    SB_LUT4 i3967_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_26_4 ), .O(n5350));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3967_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i6119_6120 (.Q(\REG.mem_63_11 ), .C(FIFO_CLK_c), .D(n6017));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10667 (.I0(rd_addr_r_c[2]), .I1(n11089), 
            .I2(n11104), .I3(rd_addr_r_c[3]), .O(n12545));
    defparam rd_addr_r_2__bdd_4_lut_10667.LUT_INIT = 16'he4aa;
    SB_LUT4 i3966_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_26_3 ), .O(n5349));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3966_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i6116_6117 (.Q(\REG.mem_63_10 ), .C(FIFO_CLK_c), .D(n6016));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6113_6114 (.Q(\REG.mem_63_9 ), .C(FIFO_CLK_c), .D(n6015));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6110_6111 (.Q(\REG.mem_63_8 ), .C(FIFO_CLK_c), .D(n6014));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6107_6108 (.Q(\REG.mem_63_7 ), .C(FIFO_CLK_c), .D(n6013));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6104_6105 (.Q(\REG.mem_63_6 ), .C(FIFO_CLK_c), .D(n6012));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6101_6102 (.Q(\REG.mem_63_5 ), .C(FIFO_CLK_c), .D(n6011));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6098_6099 (.Q(\REG.mem_63_4 ), .C(FIFO_CLK_c), .D(n6010));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6095_6096 (.Q(\REG.mem_63_3 ), .C(FIFO_CLK_c), .D(n6009));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6092_6093 (.Q(\REG.mem_63_2 ), .C(FIFO_CLK_c), .D(n6008));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6089_6090 (.Q(\REG.mem_63_1 ), .C(FIFO_CLK_c), .D(n6007));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6086_6087 (.Q(\REG.mem_63_0 ), .C(FIFO_CLK_c), .D(n6006));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6035_6036 (.Q(\REG.mem_62_15 ), .C(FIFO_CLK_c), .D(n6005));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6032_6033 (.Q(\REG.mem_62_14 ), .C(FIFO_CLK_c), .D(n6004));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6029_6030 (.Q(\REG.mem_62_13 ), .C(FIFO_CLK_c), .D(n6003));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6026_6027 (.Q(\REG.mem_62_12 ), .C(FIFO_CLK_c), .D(n6002));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i65_66 (.Q(\REG.mem_0_9 ), .C(FIFO_CLK_c), .D(n4930));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13175_bdd_4_lut (.I0(n13175), .I1(\REG.mem_25_6 ), .I2(\REG.mem_24_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11272));
    defparam n13175_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12395_bdd_4_lut (.I0(n12395), .I1(\REG.mem_37_13 ), .I2(\REG.mem_36_13 ), 
            .I3(rd_addr_r_c[1]), .O(n12398));
    defparam n12395_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12545_bdd_4_lut (.I0(n12545), .I1(n11086), .I2(n11080), .I3(rd_addr_r_c[3]), 
            .O(n11146));
    defparam n12545_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3965_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_26_2 ), .O(n5348));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3965_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9399_3_lut (.I0(\REG.mem_56_4 ), .I1(\REG.mem_57_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11237));
    defparam i9399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10687 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_7 ), 
            .I2(\REG.mem_19_7 ), .I3(rd_addr_r_c[1]), .O(n12539));
    defparam rd_addr_r_0__bdd_4_lut_10687.LUT_INIT = 16'he4aa;
    SB_LUT4 n12539_bdd_4_lut (.I0(n12539), .I1(\REG.mem_17_7 ), .I2(\REG.mem_16_7 ), 
            .I3(rd_addr_r_c[1]), .O(n12542));
    defparam n12539_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9400_3_lut (.I0(\REG.mem_58_4 ), .I1(\REG.mem_59_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11238));
    defparam i9400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10662 (.I0(rd_addr_r_c[2]), .I1(n11593), 
            .I2(n11614), .I3(rd_addr_r_c[3]), .O(n12533));
    defparam rd_addr_r_2__bdd_4_lut_10662.LUT_INIT = 16'he4aa;
    SB_DFF i68_69 (.Q(\REG.mem_0_10 ), .C(FIFO_CLK_c), .D(n4929));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i71_72 (.Q(\REG.mem_0_11 ), .C(FIFO_CLK_c), .D(n4928));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12533_bdd_4_lut (.I0(n12533), .I1(n11545), .I2(n11530), .I3(rd_addr_r_c[3]), 
            .O(n11785));
    defparam n12533_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i6023_6024 (.Q(\REG.mem_62_11 ), .C(FIFO_CLK_c), .D(n6001));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6020_6021 (.Q(\REG.mem_62_10 ), .C(FIFO_CLK_c), .D(n6000));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6017_6018 (.Q(\REG.mem_62_9 ), .C(FIFO_CLK_c), .D(n5999));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6014_6015 (.Q(\REG.mem_62_8 ), .C(FIFO_CLK_c), .D(n5998));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6011_6012 (.Q(\REG.mem_62_7 ), .C(FIFO_CLK_c), .D(n5997));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6008_6009 (.Q(\REG.mem_62_6 ), .C(FIFO_CLK_c), .D(n5996));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6005_6006 (.Q(\REG.mem_62_5 ), .C(FIFO_CLK_c), .D(n5995));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6002_6003 (.Q(\REG.mem_62_4 ), .C(FIFO_CLK_c), .D(n5994));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5999_6000 (.Q(\REG.mem_62_3 ), .C(FIFO_CLK_c), .D(n5993));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5996_5997 (.Q(\REG.mem_62_2 ), .C(FIFO_CLK_c), .D(n5992));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5993_5994 (.Q(\REG.mem_62_1 ), .C(FIFO_CLK_c), .D(n5991));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5990_5991 (.Q(\REG.mem_62_0 ), .C(FIFO_CLK_c), .D(n5990));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5939_5940 (.Q(\REG.mem_61_15 ), .C(FIFO_CLK_c), .D(n5986));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5936_5937 (.Q(\REG.mem_61_14 ), .C(FIFO_CLK_c), .D(n5985));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3964_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_26_1 ), .O(n5347));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3964_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10657 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_15 ), 
            .I2(\REG.mem_39_15 ), .I3(rd_addr_r_c[1]), .O(n12527));
    defparam rd_addr_r_0__bdd_4_lut_10657.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11185 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_11 ), 
            .I2(\REG.mem_23_11 ), .I3(rd_addr_r_c[1]), .O(n13169));
    defparam rd_addr_r_0__bdd_4_lut_11185.LUT_INIT = 16'he4aa;
    SB_LUT4 n12527_bdd_4_lut (.I0(n12527), .I1(\REG.mem_37_15 ), .I2(\REG.mem_36_15 ), 
            .I3(rd_addr_r_c[1]), .O(n12530));
    defparam n12527_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3963_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_26_0 ), .O(n5346));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3963_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13169_bdd_4_lut (.I0(n13169), .I1(\REG.mem_21_11 ), .I2(\REG.mem_20_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11653));
    defparam n13169_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10652 (.I0(rd_addr_r_c[2]), .I1(n11125), 
            .I2(n11128), .I3(rd_addr_r_c[3]), .O(n12521));
    defparam rd_addr_r_2__bdd_4_lut_10652.LUT_INIT = 16'he4aa;
    SB_LUT4 n12521_bdd_4_lut (.I0(n12521), .I1(n11119), .I2(n11113), .I3(rd_addr_r_c[3]), 
            .O(n11149));
    defparam n12521_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_11495 (.I0(rd_addr_r_c[4]), .I1(n11146), 
            .I2(n11149), .I3(rd_addr_r_c[5]), .O(n12515));
    defparam rd_addr_r_4__bdd_4_lut_11495.LUT_INIT = 16'he4aa;
    SB_LUT4 n12515_bdd_4_lut (.I0(n12515), .I1(n11137), .I2(n11131), .I3(rd_addr_r_c[5]), 
            .O(\REG.out_raw_31__N_559 [3]));
    defparam n12515_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i5933_5934 (.Q(\REG.mem_61_13 ), .C(FIFO_CLK_c), .D(n5984));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5930_5931 (.Q(\REG.mem_61_12 ), .C(FIFO_CLK_c), .D(n5983));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5927_5928 (.Q(\REG.mem_61_11 ), .C(FIFO_CLK_c), .D(n5982));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5924_5925 (.Q(\REG.mem_61_10 ), .C(FIFO_CLK_c), .D(n5981));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5921_5922 (.Q(\REG.mem_61_9 ), .C(FIFO_CLK_c), .D(n5980));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5918_5919 (.Q(\REG.mem_61_8 ), .C(FIFO_CLK_c), .D(n5979));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5915_5916 (.Q(\REG.mem_61_7 ), .C(FIFO_CLK_c), .D(n5978));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5912_5913 (.Q(\REG.mem_61_6 ), .C(FIFO_CLK_c), .D(n5977));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5909_5910 (.Q(\REG.mem_61_5 ), .C(FIFO_CLK_c), .D(n5976));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5906_5907 (.Q(\REG.mem_61_4 ), .C(FIFO_CLK_c), .D(n5975));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5903_5904 (.Q(\REG.mem_61_3 ), .C(FIFO_CLK_c), .D(n5974));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5900_5901 (.Q(\REG.mem_61_2 ), .C(FIFO_CLK_c), .D(n5973));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5897_5898 (.Q(\REG.mem_61_1 ), .C(FIFO_CLK_c), .D(n5972));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5894_5895 (.Q(\REG.mem_61_0 ), .C(FIFO_CLK_c), .D(n5971));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5843_5844 (.Q(\REG.mem_60_15 ), .C(FIFO_CLK_c), .D(n5969));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11180 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_11 ), 
            .I2(\REG.mem_27_11 ), .I3(rd_addr_r_c[1]), .O(n13163));
    defparam rd_addr_r_0__bdd_4_lut_11180.LUT_INIT = 16'he4aa;
    SB_LUT4 n13163_bdd_4_lut (.I0(n13163), .I1(\REG.mem_25_11 ), .I2(\REG.mem_24_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11656));
    defparam n13163_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3994_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_27_15 ), .O(n5377));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3994_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3993_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_27_14 ), .O(n5376));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3993_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10647 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_12 ), 
            .I2(\REG.mem_59_12 ), .I3(rd_addr_r_c[1]), .O(n12509));
    defparam rd_addr_r_0__bdd_4_lut_10647.LUT_INIT = 16'he4aa;
    SB_LUT4 i9403_3_lut (.I0(\REG.mem_62_4 ), .I1(\REG.mem_63_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11241));
    defparam i9403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9402_3_lut (.I0(\REG.mem_60_4 ), .I1(\REG.mem_61_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11240));
    defparam i9402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11275 (.I0(rd_addr_r_c[3]), .I1(n12878), 
            .I2(n11262), .I3(rd_addr_r_c[4]), .O(n13157));
    defparam rd_addr_r_3__bdd_4_lut_11275.LUT_INIT = 16'he4aa;
    SB_LUT4 n12509_bdd_4_lut (.I0(n12509), .I1(\REG.mem_57_12 ), .I2(\REG.mem_56_12 ), 
            .I3(rd_addr_r_c[1]), .O(n12512));
    defparam n12509_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3992_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_27_13 ), .O(n5375));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3992_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9821_3_lut (.I0(n13142), .I1(n13148), .I2(rd_addr_r_c[3]), 
            .I3(GND_net), .O(n11659));
    defparam i9821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13157_bdd_4_lut (.I0(n13157), .I1(n11259), .I2(n12872), .I3(rd_addr_r_c[4]), 
            .O(n13160));
    defparam n13157_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i5840_5841 (.Q(\REG.mem_60_14 ), .C(FIFO_CLK_c), .D(n5968));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10152_3_lut (.I0(\REG.mem_40_14 ), .I1(\REG.mem_41_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11990));
    defparam i10152_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5837_5838 (.Q(\REG.mem_60_13 ), .C(FIFO_CLK_c), .D(n5967));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5834_5835 (.Q(\REG.mem_60_12 ), .C(FIFO_CLK_c), .D(n5966));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5831_5832 (.Q(\REG.mem_60_11 ), .C(FIFO_CLK_c), .D(n5965));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5828_5829 (.Q(\REG.mem_60_10 ), .C(FIFO_CLK_c), .D(n5964));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5825_5826 (.Q(\REG.mem_60_9 ), .C(FIFO_CLK_c), .D(n5963));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5822_5823 (.Q(\REG.mem_60_8 ), .C(FIFO_CLK_c), .D(n5962));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5819_5820 (.Q(\REG.mem_60_7 ), .C(FIFO_CLK_c), .D(n5961));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5816_5817 (.Q(\REG.mem_60_6 ), .C(FIFO_CLK_c), .D(n5960));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5813_5814 (.Q(\REG.mem_60_5 ), .C(FIFO_CLK_c), .D(n5959));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5810_5811 (.Q(\REG.mem_60_4 ), .C(FIFO_CLK_c), .D(n5958));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5807_5808 (.Q(\REG.mem_60_3 ), .C(FIFO_CLK_c), .D(n5957));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5804_5805 (.Q(\REG.mem_60_2 ), .C(FIFO_CLK_c), .D(n5956));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5801_5802 (.Q(\REG.mem_60_1 ), .C(FIFO_CLK_c), .D(n5955));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5798_5799 (.Q(\REG.mem_60_0 ), .C(FIFO_CLK_c), .D(n5954));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync1_r__i1 (.Q(rp_sync1_r[1]), .C(FIFO_CLK_c), .D(n5953));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_LUT4 i10153_3_lut (.I0(\REG.mem_42_14 ), .I1(\REG.mem_43_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11991));
    defparam i10153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10159_3_lut (.I0(\REG.mem_46_14 ), .I1(\REG.mem_47_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11997));
    defparam i10159_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF rp_sync1_r__i2 (.Q(rp_sync1_r[2]), .C(FIFO_CLK_c), .D(n5952));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i3 (.Q(rp_sync1_r[3]), .C(FIFO_CLK_c), .D(n5951));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i4 (.Q(rp_sync1_r[4]), .C(FIFO_CLK_c), .D(n5950));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i5 (.Q(rp_sync1_r[5]), .C(FIFO_CLK_c), .D(n5949));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i6 (.Q(rp_sync1_r[6]), .C(FIFO_CLK_c), .D(n5948));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i1 (.Q(rp_sync2_r[1]), .C(FIFO_CLK_c), .D(n5947));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i2 (.Q(rp_sync2_r[2]), .C(FIFO_CLK_c), .D(n5946));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i3 (.Q(rp_sync2_r[3]), .C(FIFO_CLK_c), .D(n5945));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF i5747_5748 (.Q(\REG.mem_59_15 ), .C(FIFO_CLK_c), .D(n5944));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5744_5745 (.Q(\REG.mem_59_14 ), .C(FIFO_CLK_c), .D(n5943));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5741_5742 (.Q(\REG.mem_59_13 ), .C(FIFO_CLK_c), .D(n5942));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5738_5739 (.Q(\REG.mem_59_12 ), .C(FIFO_CLK_c), .D(n5941));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5735_5736 (.Q(\REG.mem_59_11 ), .C(FIFO_CLK_c), .D(n5940));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5732_5733 (.Q(\REG.mem_59_10 ), .C(FIFO_CLK_c), .D(n5939));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5729_5730 (.Q(\REG.mem_59_9 ), .C(FIFO_CLK_c), .D(n5938));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5726_5727 (.Q(\REG.mem_59_8 ), .C(FIFO_CLK_c), .D(n5937));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10632 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_9 ), 
            .I2(\REG.mem_55_9 ), .I3(rd_addr_r_c[1]), .O(n12503));
    defparam rd_addr_r_0__bdd_4_lut_10632.LUT_INIT = 16'he4aa;
    SB_LUT4 i3991_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_27_12 ), .O(n5374));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3991_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12503_bdd_4_lut (.I0(n12503), .I1(\REG.mem_53_9 ), .I2(\REG.mem_52_9 ), 
            .I3(rd_addr_r_c[1]), .O(n12506));
    defparam n12503_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10158_3_lut (.I0(\REG.mem_44_14 ), .I1(\REG.mem_45_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11996));
    defparam i10158_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5723_5724 (.Q(\REG.mem_59_7 ), .C(FIFO_CLK_c), .D(n5936));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5720_5721 (.Q(\REG.mem_59_6 ), .C(FIFO_CLK_c), .D(n5935));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11175 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_7 ), 
            .I2(\REG.mem_11_7 ), .I3(rd_addr_r_c[1]), .O(n13151));
    defparam rd_addr_r_0__bdd_4_lut_11175.LUT_INIT = 16'he4aa;
    SB_DFF i5717_5718 (.Q(\REG.mem_59_5 ), .C(FIFO_CLK_c), .D(n5934));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5714_5715 (.Q(\REG.mem_59_4 ), .C(FIFO_CLK_c), .D(n5933));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5711_5712 (.Q(\REG.mem_59_3 ), .C(FIFO_CLK_c), .D(n5932));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5708_5709 (.Q(\REG.mem_59_2 ), .C(FIFO_CLK_c), .D(n5931));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5705_5706 (.Q(\REG.mem_59_1 ), .C(FIFO_CLK_c), .D(n5930));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5702_5703 (.Q(\REG.mem_59_0 ), .C(FIFO_CLK_c), .D(n5929));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync2_r__i4 (.Q(rp_sync2_r[4]), .C(FIFO_CLK_c), .D(n5928));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i5 (.Q(rp_sync2_r[5]), .C(FIFO_CLK_c), .D(n5927));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i6 (.Q(rp_sync2_r[6]), .C(FIFO_CLK_c), .D(n5926));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rd_addr_r__i1 (.Q(rd_addr_r_c[1]), .C(SLM_CLK_c), .D(n5925));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i2 (.Q(rd_addr_r_c[2]), .C(SLM_CLK_c), .D(n5924));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i3 (.Q(rd_addr_r_c[3]), .C(SLM_CLK_c), .D(n5923));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i4 (.Q(rd_addr_r_c[4]), .C(SLM_CLK_c), .D(n5922));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i5 (.Q(rd_addr_r_c[5]), .C(SLM_CLK_c), .D(n5921));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i6 (.Q(\rd_addr_r[6] ), .C(SLM_CLK_c), .D(n5920));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF i5651_5652 (.Q(\REG.mem_58_15 ), .C(FIFO_CLK_c), .D(n5919));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13151_bdd_4_lut (.I0(n13151), .I1(\REG.mem_9_7 ), .I2(\REG.mem_8_7 ), 
            .I3(rd_addr_r_c[1]), .O(n13154));
    defparam n13151_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i5648_5649 (.Q(\REG.mem_58_14 ), .C(FIFO_CLK_c), .D(n5918));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i74_75 (.Q(\REG.mem_0_12 ), .C(FIFO_CLK_c), .D(n4927));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_4__bdd_4_lut_10637 (.I0(rd_addr_r_c[4]), .I1(n11764), 
            .I2(n11767), .I3(rd_addr_r_c[5]), .O(n12497));
    defparam rd_addr_r_4__bdd_4_lut_10637.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11220 (.I0(rd_addr_r_c[1]), .I1(n11093), 
            .I2(n11094), .I3(rd_addr_r_c[2]), .O(n13145));
    defparam rd_addr_r_1__bdd_4_lut_11220.LUT_INIT = 16'he4aa;
    SB_LUT4 i3990_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_27_11 ), .O(n5373));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3990_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i5645_5646 (.Q(\REG.mem_58_13 ), .C(FIFO_CLK_c), .D(n5917));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5642_5643 (.Q(\REG.mem_58_12 ), .C(FIFO_CLK_c), .D(n5916));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9378_3_lut (.I0(\REG.mem_40_4 ), .I1(\REG.mem_41_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11216));
    defparam i9378_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5639_5640 (.Q(\REG.mem_58_11 ), .C(FIFO_CLK_c), .D(n5915));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5636_5637 (.Q(\REG.mem_58_10 ), .C(FIFO_CLK_c), .D(n5914));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5633_5634 (.Q(\REG.mem_58_9 ), .C(FIFO_CLK_c), .D(n5913));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5630_5631 (.Q(\REG.mem_58_8 ), .C(FIFO_CLK_c), .D(n5912));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5627_5628 (.Q(\REG.mem_58_7 ), .C(FIFO_CLK_c), .D(n5911));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5624_5625 (.Q(\REG.mem_58_6 ), .C(FIFO_CLK_c), .D(n5910));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5621_5622 (.Q(\REG.mem_58_5 ), .C(FIFO_CLK_c), .D(n5909));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5618_5619 (.Q(\REG.mem_58_4 ), .C(FIFO_CLK_c), .D(n5908));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5615_5616 (.Q(\REG.mem_58_3 ), .C(FIFO_CLK_c), .D(n5907));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5612_5613 (.Q(\REG.mem_58_2 ), .C(FIFO_CLK_c), .D(n5906));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5609_5610 (.Q(\REG.mem_58_1 ), .C(FIFO_CLK_c), .D(n5905));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5606_5607 (.Q(\REG.mem_58_0 ), .C(FIFO_CLK_c), .D(n5904));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12497_bdd_4_lut (.I0(n12497), .I1(n11755), .I2(n11743), .I3(rd_addr_r_c[5]), 
            .O(\REG.out_raw_31__N_559 [11]));
    defparam n12497_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9379_3_lut (.I0(\REG.mem_42_4 ), .I1(\REG.mem_43_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11217));
    defparam i9379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13145_bdd_4_lut (.I0(n13145), .I1(n11001), .I2(n11000), .I3(rd_addr_r_c[2]), 
            .O(n13148));
    defparam n13145_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9382_3_lut (.I0(\REG.mem_46_4 ), .I1(\REG.mem_47_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11220));
    defparam i9382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9381_3_lut (.I0(\REG.mem_44_4 ), .I1(\REG.mem_45_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11219));
    defparam i9381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3989_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_27_10 ), .O(n5372));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3989_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9166_3_lut (.I0(n12686), .I1(n12296), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11004));
    defparam i9166_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5555_5556 (.Q(\REG.mem_57_15 ), .C(FIFO_CLK_c), .D(n5901));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5552_5553 (.Q(\REG.mem_57_14 ), .C(FIFO_CLK_c), .D(n5900));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5549_5550 (.Q(\REG.mem_57_13 ), .C(FIFO_CLK_c), .D(n5899));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5546_5547 (.Q(\REG.mem_57_12 ), .C(FIFO_CLK_c), .D(n5898));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5543_5544 (.Q(\REG.mem_57_11 ), .C(FIFO_CLK_c), .D(n5897));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5540_5541 (.Q(\REG.mem_57_10 ), .C(FIFO_CLK_c), .D(n5896));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5537_5538 (.Q(\REG.mem_57_9 ), .C(FIFO_CLK_c), .D(n5895));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5534_5535 (.Q(\REG.mem_57_8 ), .C(FIFO_CLK_c), .D(n5894));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5531_5532 (.Q(\REG.mem_57_7 ), .C(FIFO_CLK_c), .D(n5893));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5528_5529 (.Q(\REG.mem_57_6 ), .C(FIFO_CLK_c), .D(n5892));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5525_5526 (.Q(\REG.mem_57_5 ), .C(FIFO_CLK_c), .D(n5891));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5522_5523 (.Q(\REG.mem_57_4 ), .C(FIFO_CLK_c), .D(n5890));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5519_5520 (.Q(\REG.mem_57_3 ), .C(FIFO_CLK_c), .D(n5889));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5516_5517 (.Q(\REG.mem_57_2 ), .C(FIFO_CLK_c), .D(n5888));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5513_5514 (.Q(\REG.mem_57_1 ), .C(FIFO_CLK_c), .D(n5887));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut (.I0(rd_addr_r[0]), .I1(\REG.mem_18_1 ), 
            .I2(\REG.mem_19_1 ), .I3(rd_addr_r_c[1]), .O(n13859));
    defparam rd_addr_r_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n13859_bdd_4_lut (.I0(n13859), .I1(\REG.mem_17_1 ), .I2(\REG.mem_16_1 ), 
            .I3(rd_addr_r_c[1]), .O(n11389));
    defparam n13859_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3988_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_27_9 ), .O(n5371));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3988_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11160 (.I0(rd_addr_r_c[1]), .I1(n12023), 
            .I2(n12024), .I3(rd_addr_r_c[2]), .O(n13139));
    defparam rd_addr_r_1__bdd_4_lut_11160.LUT_INIT = 16'he4aa;
    SB_DFF i5510_5511 (.Q(\REG.mem_57_0 ), .C(FIFO_CLK_c), .D(n5885));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3987_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_27_8 ), .O(n5370));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3987_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i5459_5460 (.Q(\REG.mem_56_15 ), .C(FIFO_CLK_c), .D(n5884));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5456_5457 (.Q(\REG.mem_56_14 ), .C(FIFO_CLK_c), .D(n5883));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5453_5454 (.Q(\REG.mem_56_13 ), .C(FIFO_CLK_c), .D(n5882));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5450_5451 (.Q(\REG.mem_56_12 ), .C(FIFO_CLK_c), .D(n5881));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5447_5448 (.Q(\REG.mem_56_11 ), .C(FIFO_CLK_c), .D(n5880));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5444_5445 (.Q(\REG.mem_56_10 ), .C(FIFO_CLK_c), .D(n5879));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5441_5442 (.Q(\REG.mem_56_9 ), .C(FIFO_CLK_c), .D(n5878));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5438_5439 (.Q(\REG.mem_56_8 ), .C(FIFO_CLK_c), .D(n5877));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5435_5436 (.Q(\REG.mem_56_7 ), .C(FIFO_CLK_c), .D(n5876));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5432_5433 (.Q(\REG.mem_56_6 ), .C(FIFO_CLK_c), .D(n5875));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5429_5430 (.Q(\REG.mem_56_5 ), .C(FIFO_CLK_c), .D(n5874));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5426_5427 (.Q(\REG.mem_56_4 ), .C(FIFO_CLK_c), .D(n5873));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5423_5424 (.Q(\REG.mem_56_3 ), .C(FIFO_CLK_c), .D(n5872));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5420_5421 (.Q(\REG.mem_56_2 ), .C(FIFO_CLK_c), .D(n5871));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5417_5418 (.Q(\REG.mem_56_1 ), .C(FIFO_CLK_c), .D(n5870));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9798_3_lut (.I0(\REG.mem_32_8 ), .I1(\REG.mem_33_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11636));
    defparam i9798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9799_3_lut (.I0(\REG.mem_34_8 ), .I1(\REG.mem_35_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11637));
    defparam i9799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13139_bdd_4_lut (.I0(n13139), .I1(n12012), .I2(n12011), .I3(rd_addr_r_c[2]), 
            .O(n13142));
    defparam n13139_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9844_3_lut (.I0(\REG.mem_38_8 ), .I1(\REG.mem_39_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11682));
    defparam i9844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11755 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_14 ), 
            .I2(\REG.mem_59_14 ), .I3(rd_addr_r_c[1]), .O(n13853));
    defparam rd_addr_r_0__bdd_4_lut_11755.LUT_INIT = 16'he4aa;
    SB_LUT4 i9843_3_lut (.I0(\REG.mem_36_8 ), .I1(\REG.mem_37_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11681));
    defparam i9843_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5414_5415 (.Q(\REG.mem_56_0 ), .C(FIFO_CLK_c), .D(n5865));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wp_sync1_r__i1 (.Q(wp_sync1_r[1]), .C(SLM_CLK_c), .D(n5864));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i2 (.Q(wp_sync1_r[2]), .C(SLM_CLK_c), .D(n5863));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i3 (.Q(wp_sync1_r[3]), .C(SLM_CLK_c), .D(n5862));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i4 (.Q(wp_sync1_r[4]), .C(SLM_CLK_c), .D(n5861));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i5 (.Q(wp_sync1_r[5]), .C(SLM_CLK_c), .D(n5860));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i6 (.Q(wp_sync1_r[6]), .C(SLM_CLK_c), .D(n5859));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF i5363_5364 (.Q(\REG.mem_55_15 ), .C(FIFO_CLK_c), .D(n5858));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5360_5361 (.Q(\REG.mem_55_14 ), .C(FIFO_CLK_c), .D(n5857));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5357_5358 (.Q(\REG.mem_55_13 ), .C(FIFO_CLK_c), .D(n5856));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5354_5355 (.Q(\REG.mem_55_12 ), .C(FIFO_CLK_c), .D(n5855));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5351_5352 (.Q(\REG.mem_55_11 ), .C(FIFO_CLK_c), .D(n5854));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5348_5349 (.Q(\REG.mem_55_10 ), .C(FIFO_CLK_c), .D(n5853));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY wr_addr_r_6__I_0_141_7 (.CI(n10137), .I0(wr_addr_r[5]), .I1(GND_net), 
            .CO(n10138));
    SB_LUT4 wr_addr_r_6__I_0_141_6_lut (.I0(GND_net), .I1(wr_addr_r[4]), 
            .I2(GND_net), .I3(n10136), .O(wr_addr_p1_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_141_6 (.CI(n10136), .I0(wr_addr_r[4]), .I1(GND_net), 
            .CO(n10137));
    SB_LUT4 wr_addr_r_6__I_0_141_5_lut (.I0(GND_net), .I1(wr_addr_r[3]), 
            .I2(GND_net), .I3(n10135), .O(wr_addr_p1_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_141_5 (.CI(n10135), .I0(wr_addr_r[3]), .I1(GND_net), 
            .CO(n10136));
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_3 (.CI(n10090), .I0(wp_sync_w[1]), 
            .I1(n1[1]), .CO(n10091));
    SB_LUT4 wr_addr_r_6__I_0_141_4_lut (.I0(GND_net), .I1(wr_addr_r[2]), 
            .I2(GND_net), .I3(n10134), .O(wr_addr_p1_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_2_lut (.I0(GND_net), .I1(wp_sync_w[0]), 
            .I2(n1[0]), .I3(VCC_net), .O(\rd_sig_diff0_w[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_141_4 (.CI(n10134), .I0(wr_addr_r[2]), .I1(GND_net), 
            .CO(n10135));
    SB_DFF i5345_5346 (.Q(\REG.mem_55_9 ), .C(FIFO_CLK_c), .D(n5852));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5342_5343 (.Q(\REG.mem_55_8 ), .C(FIFO_CLK_c), .D(n5851));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5339_5340 (.Q(\REG.mem_55_7 ), .C(FIFO_CLK_c), .D(n5850));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5336_5337 (.Q(\REG.mem_55_6 ), .C(FIFO_CLK_c), .D(n5849));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5333_5334 (.Q(\REG.mem_55_5 ), .C(FIFO_CLK_c), .D(n5848));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5330_5331 (.Q(\REG.mem_55_4 ), .C(FIFO_CLK_c), .D(n5847));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5327_5328 (.Q(\REG.mem_55_3 ), .C(FIFO_CLK_c), .D(n5846));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5324_5325 (.Q(\REG.mem_55_2 ), .C(FIFO_CLK_c), .D(n5845));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5321_5322 (.Q(\REG.mem_55_1 ), .C(FIFO_CLK_c), .D(n5844));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5318_5319 (.Q(\REG.mem_55_0 ), .C(FIFO_CLK_c), .D(n5843));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wp_sync2_r__i1 (.Q(wp_sync2_r[1]), .C(SLM_CLK_c), .D(n5842));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i2 (.Q(wp_sync2_r[2]), .C(SLM_CLK_c), .D(n5841));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i3 (.Q(wp_sync2_r[3]), .C(SLM_CLK_c), .D(n5839));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i4 (.Q(wp_sync2_r[4]), .C(SLM_CLK_c), .D(n5838));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i5 (.Q(wp_sync2_r[5]), .C(SLM_CLK_c), .D(n5837));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_LUT4 wr_addr_r_6__I_0_141_3_lut (.I0(GND_net), .I1(wr_addr_r[1]), 
            .I2(GND_net), .I3(n10133), .O(wr_addr_p1_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_r_6__I_0_151_8_lut (.I0(GND_net), .I1(\rd_addr_r[6] ), 
            .I2(GND_net), .I3(n10144), .O(rd_addr_p1_w[6])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_141_3 (.CI(n10133), .I0(wr_addr_r[1]), .I1(GND_net), 
            .CO(n10134));
    SB_LUT4 wr_addr_r_6__I_0_141_2_lut (.I0(GND_net), .I1(wr_addr_r[0]), 
            .I2(GND_net), .I3(VCC_net), .O(wr_addr_p1_w[0])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_r_6__I_0_151_7_lut (.I0(GND_net), .I1(rd_addr_r_c[5]), 
            .I2(GND_net), .I3(n10143), .O(rd_addr_p1_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_141_2 (.CI(VCC_net), .I0(wr_addr_r[0]), .I1(GND_net), 
            .CO(n10133));
    SB_LUT4 i9855_3_lut (.I0(\REG.mem_16_15 ), .I1(\REG.mem_17_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11693));
    defparam i9855_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rd_addr_r_6__I_0_151_7 (.CI(n10143), .I0(rd_addr_r_c[5]), .I1(GND_net), 
            .CO(n10144));
    SB_LUT4 i9856_3_lut (.I0(\REG.mem_18_15 ), .I1(\REG.mem_19_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11694));
    defparam i9856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_add_2_8_lut (.I0(n10979), .I1(wr_grey_sync_r[6]), 
            .I2(n1_adj_45[6]), .I3(n10101), .O(\afull_flag_impl.af_flag_nxt_w )) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i9877_3_lut (.I0(\REG.mem_22_15 ), .I1(\REG.mem_23_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11715));
    defparam i9877_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF wp_sync2_r__i6 (.Q(wp_sync2_r[6]), .C(SLM_CLK_c), .D(n5836));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF i5267_5268 (.Q(\REG.mem_54_15 ), .C(FIFO_CLK_c), .D(n5835));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5264_5265 (.Q(\REG.mem_54_14 ), .C(FIFO_CLK_c), .D(n5834));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5261_5262 (.Q(\REG.mem_54_13 ), .C(FIFO_CLK_c), .D(n5833));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5258_5259 (.Q(\REG.mem_54_12 ), .C(FIFO_CLK_c), .D(n5832));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5255_5256 (.Q(\REG.mem_54_11 ), .C(FIFO_CLK_c), .D(n5831));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5252_5253 (.Q(\REG.mem_54_10 ), .C(FIFO_CLK_c), .D(n5830));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5249_5250 (.Q(\REG.mem_54_9 ), .C(FIFO_CLK_c), .D(n5829));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5246_5247 (.Q(\REG.mem_54_8 ), .C(FIFO_CLK_c), .D(n5828));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5243_5244 (.Q(\REG.mem_54_7 ), .C(FIFO_CLK_c), .D(n5827));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5240_5241 (.Q(\REG.mem_54_6 ), .C(FIFO_CLK_c), .D(n5826));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5237_5238 (.Q(\REG.mem_54_5 ), .C(FIFO_CLK_c), .D(n5825));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5234_5235 (.Q(\REG.mem_54_4 ), .C(FIFO_CLK_c), .D(n5824));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5231_5232 (.Q(\REG.mem_54_3 ), .C(FIFO_CLK_c), .D(n5823));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5228_5229 (.Q(\REG.mem_54_2 ), .C(FIFO_CLK_c), .D(n5822));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5225_5226 (.Q(\REG.mem_54_1 ), .C(FIFO_CLK_c), .D(n5821));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9876_3_lut (.I0(\REG.mem_20_15 ), .I1(\REG.mem_21_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11714));
    defparam i9876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_add_2_7_lut (.I0(n10951), .I1(wr_addr_r[5]), 
            .I2(rp_sync_w[5]), .I3(n10100), .O(n10979)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY wr_addr_r_6__I_0_add_2_7 (.CI(n10100), .I0(wr_addr_r[5]), .I1(rp_sync_w[5]), 
            .CO(n10101));
    SB_LUT4 rd_addr_r_6__I_0_151_6_lut (.I0(GND_net), .I1(rd_addr_r_c[4]), 
            .I2(GND_net), .I3(n10142), .O(rd_addr_p1_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wr_addr_r_6__I_0_add_2_6_lut (.I0(n2_adj_22), .I1(wr_addr_r[4]), 
            .I2(rp_sync_w[4]), .I3(n10099), .O(n10925)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_6_lut.LUT_INIT = 16'hebbe;
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_2 (.CI(VCC_net), .I0(wp_sync_w[0]), 
            .I1(n1[0]), .CO(n10090));
    SB_CARRY wr_addr_r_6__I_0_add_2_6 (.CI(n10099), .I0(wr_addr_r[4]), .I1(rp_sync_w[4]), 
            .CO(n10100));
    SB_LUT4 i9354_3_lut (.I0(\REG.mem_24_4 ), .I1(\REG.mem_25_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11192));
    defparam i9354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_add_2_5_lut (.I0(GND_net), .I1(wr_addr_r[3]), 
            .I2(rp_sync_w[3]), .I3(n10098), .O(wr_sig_diff0_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_add_2_5 (.CI(n10098), .I0(wr_addr_r[3]), .I1(rp_sync_w[3]), 
            .CO(n10099));
    SB_LUT4 i9355_3_lut (.I0(\REG.mem_26_4 ), .I1(\REG.mem_27_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11193));
    defparam i9355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10068_3_lut (.I0(\REG.mem_32_2 ), .I1(\REG.mem_33_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11906));
    defparam i10068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10069_3_lut (.I0(\REG.mem_34_2 ), .I1(\REG.mem_35_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11907));
    defparam i10069_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rd_addr_r_6__I_0_151_6 (.CI(n10142), .I0(rd_addr_r_c[4]), .I1(GND_net), 
            .CO(n10143));
    SB_LUT4 i9361_3_lut (.I0(\REG.mem_30_4 ), .I1(\REG.mem_31_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11199));
    defparam i9361_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5222_5223 (.Q(\REG.mem_54_0 ), .C(FIFO_CLK_c), .D(n5820));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5171_5172 (.Q(\REG.mem_53_15 ), .C(FIFO_CLK_c), .D(n5819));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5168_5169 (.Q(\REG.mem_53_14 ), .C(FIFO_CLK_c), .D(n5818));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5165_5166 (.Q(\REG.mem_53_13 ), .C(FIFO_CLK_c), .D(n5817));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5162_5163 (.Q(\REG.mem_53_12 ), .C(FIFO_CLK_c), .D(n5816));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5159_5160 (.Q(\REG.mem_53_11 ), .C(FIFO_CLK_c), .D(n5815));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5156_5157 (.Q(\REG.mem_53_10 ), .C(FIFO_CLK_c), .D(n5814));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5153_5154 (.Q(\REG.mem_53_9 ), .C(FIFO_CLK_c), .D(n5813));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5150_5151 (.Q(\REG.mem_53_8 ), .C(FIFO_CLK_c), .D(n5812));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5147_5148 (.Q(\REG.mem_53_7 ), .C(FIFO_CLK_c), .D(n5811));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5144_5145 (.Q(\REG.mem_53_6 ), .C(FIFO_CLK_c), .D(n5810));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5141_5142 (.Q(\REG.mem_53_5 ), .C(FIFO_CLK_c), .D(n5809));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5138_5139 (.Q(\REG.mem_53_4 ), .C(FIFO_CLK_c), .D(n5808));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5135_5136 (.Q(\REG.mem_53_3 ), .C(FIFO_CLK_c), .D(n5807));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5132_5133 (.Q(\REG.mem_53_2 ), .C(FIFO_CLK_c), .D(n5806));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5129_5130 (.Q(\REG.mem_53_1 ), .C(FIFO_CLK_c), .D(n5805));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9360_3_lut (.I0(\REG.mem_28_4 ), .I1(\REG.mem_29_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11198));
    defparam i9360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10072_3_lut (.I0(\REG.mem_38_2 ), .I1(\REG.mem_39_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11910));
    defparam i10072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_6__I_0_151_5_lut (.I0(GND_net), .I1(rd_addr_r_c[3]), 
            .I2(GND_net), .I3(n10141), .O(rd_addr_p1_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10071_3_lut (.I0(\REG.mem_36_2 ), .I1(\REG.mem_37_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11909));
    defparam i10071_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rd_addr_r_6__I_0_151_5 (.CI(n10141), .I0(rd_addr_r_c[3]), .I1(GND_net), 
            .CO(n10142));
    SB_DFF i5126_5127 (.Q(\REG.mem_53_0 ), .C(FIFO_CLK_c), .D(n5804));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5075_5076 (.Q(\REG.mem_52_15 ), .C(FIFO_CLK_c), .D(n5803));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5072_5073 (.Q(\REG.mem_52_14 ), .C(FIFO_CLK_c), .D(n5802));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5069_5070 (.Q(\REG.mem_52_13 ), .C(FIFO_CLK_c), .D(n5801));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5066_5067 (.Q(\REG.mem_52_12 ), .C(FIFO_CLK_c), .D(n5800));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5063_5064 (.Q(\REG.mem_52_11 ), .C(FIFO_CLK_c), .D(n5799));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5060_5061 (.Q(\REG.mem_52_10 ), .C(FIFO_CLK_c), .D(n5798));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5057_5058 (.Q(\REG.mem_52_9 ), .C(FIFO_CLK_c), .D(n5797));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5054_5055 (.Q(\REG.mem_52_8 ), .C(FIFO_CLK_c), .D(n5796));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5051_5052 (.Q(\REG.mem_52_7 ), .C(FIFO_CLK_c), .D(n5795));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5048_5049 (.Q(\REG.mem_52_6 ), .C(FIFO_CLK_c), .D(n5794));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5045_5046 (.Q(\REG.mem_52_5 ), .C(FIFO_CLK_c), .D(n5793));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5042_5043 (.Q(\REG.mem_52_4 ), .C(FIFO_CLK_c), .D(n5792));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5039_5040 (.Q(\REG.mem_52_3 ), .C(FIFO_CLK_c), .D(n5791));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5036_5037 (.Q(\REG.mem_52_2 ), .C(FIFO_CLK_c), .D(n5790));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5033_5034 (.Q(\REG.mem_52_1 ), .C(FIFO_CLK_c), .D(n5789));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11165 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_15 ), 
            .I2(\REG.mem_11_15 ), .I3(rd_addr_r_c[1]), .O(n13133));
    defparam rd_addr_r_0__bdd_4_lut_11165.LUT_INIT = 16'he4aa;
    SB_LUT4 i10104_3_lut (.I0(\REG.mem_48_2 ), .I1(\REG.mem_49_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11942));
    defparam i10104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3986_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_27_7 ), .O(n5369));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3986_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10105_3_lut (.I0(\REG.mem_50_2 ), .I1(\REG.mem_51_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11943));
    defparam i10105_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13853_bdd_4_lut (.I0(n13853), .I1(\REG.mem_57_14 ), .I2(\REG.mem_56_14 ), 
            .I3(rd_addr_r_c[1]), .O(n10993));
    defparam n13853_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10111_3_lut (.I0(\REG.mem_54_2 ), .I1(\REG.mem_55_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11949));
    defparam i10111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_add_2_4_lut (.I0(GND_net), .I1(wr_addr_r[2]), 
            .I2(rp_sync_w[2]), .I3(n10097), .O(wr_sig_diff0_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF i5030_5031 (.Q(\REG.mem_52_0 ), .C(FIFO_CLK_c), .D(n5788));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY wr_addr_r_6__I_0_add_2_4 (.CI(n10097), .I0(wr_addr_r[2]), .I1(rp_sync_w[2]), 
            .CO(n10098));
    SB_DFF i4979_4980 (.Q(\REG.mem_51_15 ), .C(FIFO_CLK_c), .D(n5787));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4976_4977 (.Q(\REG.mem_51_14 ), .C(FIFO_CLK_c), .D(n5786));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4973_4974 (.Q(\REG.mem_51_13 ), .C(FIFO_CLK_c), .D(n5785));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4970_4971 (.Q(\REG.mem_51_12 ), .C(FIFO_CLK_c), .D(n5784));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4967_4968 (.Q(\REG.mem_51_11 ), .C(FIFO_CLK_c), .D(n5783));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4964_4965 (.Q(\REG.mem_51_10 ), .C(FIFO_CLK_c), .D(n5782));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4961_4962 (.Q(\REG.mem_51_9 ), .C(FIFO_CLK_c), .D(n5781));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4958_4959 (.Q(\REG.mem_51_8 ), .C(FIFO_CLK_c), .D(n5780));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4955_4956 (.Q(\REG.mem_51_7 ), .C(FIFO_CLK_c), .D(n5779));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4952_4953 (.Q(\REG.mem_51_6 ), .C(FIFO_CLK_c), .D(n5778));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4949_4950 (.Q(\REG.mem_51_5 ), .C(FIFO_CLK_c), .D(n5777));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4946_4947 (.Q(\REG.mem_51_4 ), .C(FIFO_CLK_c), .D(n5776));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4943_4944 (.Q(\REG.mem_51_3 ), .C(FIFO_CLK_c), .D(n5775));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4940_4941 (.Q(\REG.mem_51_2 ), .C(FIFO_CLK_c), .D(n5774));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4937_4938 (.Q(\REG.mem_51_1 ), .C(FIFO_CLK_c), .D(n5773));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10110_3_lut (.I0(\REG.mem_52_2 ), .I1(\REG.mem_53_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11948));
    defparam i10110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_add_2_3_lut (.I0(GND_net), .I1(wr_addr_r[1]), 
            .I2(rp_sync_w[1]), .I3(n10096), .O(wr_sig_diff0_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_add_2_3 (.CI(n10096), .I0(wr_addr_r[1]), .I1(rp_sync_w[1]), 
            .CO(n10097));
    SB_LUT4 i9330_3_lut (.I0(\REG.mem_8_4 ), .I1(\REG.mem_9_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11168));
    defparam i9330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9331_3_lut (.I0(\REG.mem_10_4 ), .I1(\REG.mem_11_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11169));
    defparam i9331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_6__I_0_151_4_lut (.I0(GND_net), .I1(rd_addr_r_c[2]), 
            .I2(GND_net), .I3(n10140), .O(rd_addr_p1_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wr_addr_r_6__I_0_add_2_2_lut (.I0(GND_net), .I1(wr_addr_r[0]), 
            .I2(rp_sync_w[0]), .I3(VCC_net), .O(wr_sig_diff0_w[0])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF i4934_4935 (.Q(\REG.mem_51_0 ), .C(FIFO_CLK_c), .D(n5772));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4883_4884 (.Q(\REG.mem_50_15 ), .C(FIFO_CLK_c), .D(n5771));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4880_4881 (.Q(\REG.mem_50_14 ), .C(FIFO_CLK_c), .D(n5770));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4877_4878 (.Q(\REG.mem_50_13 ), .C(FIFO_CLK_c), .D(n5769));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4874_4875 (.Q(\REG.mem_50_12 ), .C(FIFO_CLK_c), .D(n5768));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4871_4872 (.Q(\REG.mem_50_11 ), .C(FIFO_CLK_c), .D(n5767));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4868_4869 (.Q(\REG.mem_50_10 ), .C(FIFO_CLK_c), .D(n5766));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4865_4866 (.Q(\REG.mem_50_9 ), .C(FIFO_CLK_c), .D(n5765));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4862_4863 (.Q(\REG.mem_50_8 ), .C(FIFO_CLK_c), .D(n5764));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4859_4860 (.Q(\REG.mem_50_7 ), .C(FIFO_CLK_c), .D(n5763));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4856_4857 (.Q(\REG.mem_50_6 ), .C(FIFO_CLK_c), .D(n5762));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4853_4854 (.Q(\REG.mem_50_5 ), .C(FIFO_CLK_c), .D(n5761));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4850_4851 (.Q(\REG.mem_50_4 ), .C(FIFO_CLK_c), .D(n5760));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4847_4848 (.Q(\REG.mem_50_3 ), .C(FIFO_CLK_c), .D(n5759));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4844_4845 (.Q(\REG.mem_50_2 ), .C(FIFO_CLK_c), .D(n5758));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4841_4842 (.Q(\REG.mem_50_1 ), .C(FIFO_CLK_c), .D(n5757));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY wr_addr_r_6__I_0_add_2_2 (.CI(VCC_net), .I0(wr_addr_r[0]), 
            .I1(rp_sync_w[0]), .CO(n10096));
    SB_LUT4 i9334_3_lut (.I0(\REG.mem_14_4 ), .I1(\REG.mem_15_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11172));
    defparam i9334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_8_lut (.I0(rd_sig_diff0_w[5]), .I1(wp_sync2_r[6]), 
            .I2(n1[6]), .I3(n10095), .O(n10873)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_7_lut (.I0(GND_net), .I1(wp_sync_w[5]), 
            .I2(n1[5]), .I3(n10094), .O(rd_sig_diff0_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9333_3_lut (.I0(\REG.mem_12_4 ), .I1(\REG.mem_13_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11171));
    defparam i9333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10011_3_lut (.I0(\REG.mem_0_14 ), .I1(\REG.mem_1_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11849));
    defparam i10011_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rd_addr_r_6__I_0_151_4 (.CI(n10140), .I0(rd_addr_r_c[2]), .I1(GND_net), 
            .CO(n10141));
    SB_DFF \REG.out_buffer__i14  (.Q(\fifo_data_out[14] ), .C(SLM_CLK_c), 
           .D(n10582));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i15  (.Q(\fifo_data_out[15] ), .C(SLM_CLK_c), 
           .D(n10588));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF i4838_4839 (.Q(\REG.mem_50_0 ), .C(FIFO_CLK_c), .D(n5753));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4787_4788 (.Q(\REG.mem_49_15 ), .C(FIFO_CLK_c), .D(n5752));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4784_4785 (.Q(\REG.mem_49_14 ), .C(FIFO_CLK_c), .D(n5751));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4781_4782 (.Q(\REG.mem_49_13 ), .C(FIFO_CLK_c), .D(n5750));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4778_4779 (.Q(\REG.mem_49_12 ), .C(FIFO_CLK_c), .D(n5749));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4775_4776 (.Q(\REG.mem_49_11 ), .C(FIFO_CLK_c), .D(n5748));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4772_4773 (.Q(\REG.mem_49_10 ), .C(FIFO_CLK_c), .D(n5747));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4769_4770 (.Q(\REG.mem_49_9 ), .C(FIFO_CLK_c), .D(n5746));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4766_4767 (.Q(\REG.mem_49_8 ), .C(FIFO_CLK_c), .D(n5745));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4763_4764 (.Q(\REG.mem_49_7 ), .C(FIFO_CLK_c), .D(n5744));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4760_4761 (.Q(\REG.mem_49_6 ), .C(FIFO_CLK_c), .D(n5743));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4757_4758 (.Q(\REG.mem_49_5 ), .C(FIFO_CLK_c), .D(n5742));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4754_4755 (.Q(\REG.mem_49_4 ), .C(FIFO_CLK_c), .D(n5741));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10012_3_lut (.I0(\REG.mem_2_14 ), .I1(\REG.mem_3_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11850));
    defparam i10012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_6__I_0_151_3_lut (.I0(GND_net), .I1(rd_addr_r_c[1]), 
            .I2(GND_net), .I3(n10139), .O(rd_addr_p1_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10015_3_lut (.I0(\REG.mem_6_14 ), .I1(\REG.mem_7_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11853));
    defparam i10015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10014_3_lut (.I0(\REG.mem_4_14 ), .I1(\REG.mem_5_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11852));
    defparam i10014_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rd_addr_r_6__I_0_151_3 (.CI(n10139), .I0(rd_addr_r_c[1]), .I1(GND_net), 
            .CO(n10140));
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_7 (.CI(n10094), .I0(wp_sync_w[5]), 
            .I1(n1[5]), .CO(n10095));
    SB_DFF i4751_4752 (.Q(\REG.mem_49_3 ), .C(FIFO_CLK_c), .D(n5740));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4748_4749 (.Q(\REG.mem_49_2 ), .C(FIFO_CLK_c), .D(n5739));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4745_4746 (.Q(\REG.mem_49_1 ), .C(FIFO_CLK_c), .D(n5738));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4742_4743 (.Q(\REG.mem_49_0 ), .C(FIFO_CLK_c), .D(n5737));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4691_4692 (.Q(\REG.mem_48_15 ), .C(FIFO_CLK_c), .D(n5736));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4688_4689 (.Q(\REG.mem_48_14 ), .C(FIFO_CLK_c), .D(n5735));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4685_4686 (.Q(\REG.mem_48_13 ), .C(FIFO_CLK_c), .D(n5734));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4682_4683 (.Q(\REG.mem_48_12 ), .C(FIFO_CLK_c), .D(n5733));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4679_4680 (.Q(\REG.mem_48_11 ), .C(FIFO_CLK_c), .D(n5732));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4676_4677 (.Q(\REG.mem_48_10 ), .C(FIFO_CLK_c), .D(n5731));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4673_4674 (.Q(\REG.mem_48_9 ), .C(FIFO_CLK_c), .D(n5730));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4670_4671 (.Q(\REG.mem_48_8 ), .C(FIFO_CLK_c), .D(n5729));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4667_4668 (.Q(\REG.mem_48_7 ), .C(FIFO_CLK_c), .D(n5728));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4664_4665 (.Q(\REG.mem_48_6 ), .C(FIFO_CLK_c), .D(n5727));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4661_4662 (.Q(\REG.mem_48_5 ), .C(FIFO_CLK_c), .D(n5726));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9171_3_lut (.I0(n12446), .I1(n12386), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11009));
    defparam i9171_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i4658_4659 (.Q(\REG.mem_48_4 ), .C(FIFO_CLK_c), .D(n5725));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4655_4656 (.Q(\REG.mem_48_3 ), .C(FIFO_CLK_c), .D(n5724));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_6_lut (.I0(rd_sig_diff0_w[3]), .I1(wp_sync_w[4]), 
            .I2(n1[4]), .I3(n10093), .O(n10877)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_6_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 n13133_bdd_4_lut (.I0(n13133), .I1(\REG.mem_9_15 ), .I2(\REG.mem_8_15 ), 
            .I3(rd_addr_r_c[1]), .O(n13136));
    defparam n13133_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11750 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_7 ), 
            .I2(\REG.mem_31_7 ), .I3(rd_addr_r_c[1]), .O(n13847));
    defparam rd_addr_r_0__bdd_4_lut_11750.LUT_INIT = 16'he4aa;
    SB_DFF i4652_4653 (.Q(\REG.mem_48_2 ), .C(FIFO_CLK_c), .D(n5723));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4649_4650 (.Q(\REG.mem_48_1 ), .C(FIFO_CLK_c), .D(n5722));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4646_4647 (.Q(\REG.mem_48_0 ), .C(FIFO_CLK_c), .D(n5721));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4595_4596 (.Q(\REG.mem_47_15 ), .C(FIFO_CLK_c), .D(n5720));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13847_bdd_4_lut (.I0(n13847), .I1(\REG.mem_29_7 ), .I2(\REG.mem_28_7 ), 
            .I3(rd_addr_r_c[1]), .O(n13850));
    defparam n13847_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4592_4593 (.Q(\REG.mem_47_14 ), .C(FIFO_CLK_c), .D(n5719));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i77_78 (.Q(\REG.mem_0_13 ), .C(FIFO_CLK_c), .D(n4926));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i80_81 (.Q(\REG.mem_0_14 ), .C(FIFO_CLK_c), .D(n4925));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9172_3_lut (.I0(n12368), .I1(n12350), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11010));
    defparam i9172_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i4589_4590 (.Q(\REG.mem_47_13 ), .C(FIFO_CLK_c), .D(n5718));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4586_4587 (.Q(\REG.mem_47_12 ), .C(FIFO_CLK_c), .D(n5717));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4583_4584 (.Q(\REG.mem_47_11 ), .C(FIFO_CLK_c), .D(n5716));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4580_4581 (.Q(\REG.mem_47_10 ), .C(FIFO_CLK_c), .D(n5715));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4577_4578 (.Q(\REG.mem_47_9 ), .C(FIFO_CLK_c), .D(n5714));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4574_4575 (.Q(\REG.mem_47_8 ), .C(FIFO_CLK_c), .D(n5713));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4571_4572 (.Q(\REG.mem_47_7 ), .C(FIFO_CLK_c), .D(n5712));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4568_4569 (.Q(\REG.mem_47_6 ), .C(FIFO_CLK_c), .D(n5711));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4565_4566 (.Q(\REG.mem_47_5 ), .C(FIFO_CLK_c), .D(n5710));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4562_4563 (.Q(\REG.mem_47_4 ), .C(FIFO_CLK_c), .D(n5709));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4559_4560 (.Q(\REG.mem_47_3 ), .C(FIFO_CLK_c), .D(n5708));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4556_4557 (.Q(\REG.mem_47_2 ), .C(FIFO_CLK_c), .D(n5707));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4553_4554 (.Q(\REG.mem_47_1 ), .C(FIFO_CLK_c), .D(n5706));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4550_4551 (.Q(\REG.mem_47_0 ), .C(FIFO_CLK_c), .D(n5705));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4499_4500 (.Q(\REG.mem_46_15 ), .C(FIFO_CLK_c), .D(n5704));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4496_4497 (.Q(\REG.mem_46_14 ), .C(FIFO_CLK_c), .D(n5703));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10627 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_0 ), 
            .I2(\REG.mem_63_0 ), .I3(rd_addr_r_c[1]), .O(n12479));
    defparam rd_addr_r_0__bdd_4_lut_10627.LUT_INIT = 16'he4aa;
    SB_DFF i83_84 (.Q(\REG.mem_0_15 ), .C(FIFO_CLK_c), .D(n4924));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12479_bdd_4_lut (.I0(n12479), .I1(\REG.mem_61_0 ), .I2(\REG.mem_60_0 ), 
            .I3(rd_addr_r_c[1]), .O(n12482));
    defparam n12479_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut (.I0(rd_addr_r_c[2]), .I1(n12422), .I2(n12380), 
            .I3(rd_addr_r_c[3]), .O(n13841));
    defparam rd_addr_r_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11150 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_12 ), 
            .I2(\REG.mem_31_12 ), .I3(rd_addr_r_c[1]), .O(n13127));
    defparam rd_addr_r_0__bdd_4_lut_11150.LUT_INIT = 16'he4aa;
    SB_DFF i4493_4494 (.Q(\REG.mem_46_13 ), .C(FIFO_CLK_c), .D(n5702));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9174_3_lut (.I0(n12338), .I1(n13814), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11012));
    defparam i9174_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i4490_4491 (.Q(\REG.mem_46_12 ), .C(FIFO_CLK_c), .D(n5701));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4487_4488 (.Q(\REG.mem_46_11 ), .C(FIFO_CLK_c), .D(n5700));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13841_bdd_4_lut (.I0(n13841), .I1(n12506), .I2(n12620), .I3(rd_addr_r_c[3]), 
            .O(n11401));
    defparam n13841_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4484_4485 (.Q(\REG.mem_46_10 ), .C(FIFO_CLK_c), .D(n5699));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3985_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_27_6 ), .O(n5368));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3985_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i4481_4482 (.Q(\REG.mem_46_9 ), .C(FIFO_CLK_c), .D(n5698));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13127_bdd_4_lut (.I0(n13127), .I1(\REG.mem_29_12 ), .I2(\REG.mem_28_12 ), 
            .I3(rd_addr_r_c[1]), .O(n13130));
    defparam n13127_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4478_4479 (.Q(\REG.mem_46_8 ), .C(FIFO_CLK_c), .D(n5697));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4475_4476 (.Q(\REG.mem_46_7 ), .C(FIFO_CLK_c), .D(n5696));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4472_4473 (.Q(\REG.mem_46_6 ), .C(FIFO_CLK_c), .D(n5695));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11145 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_3 ), 
            .I2(\REG.mem_55_3 ), .I3(rd_addr_r_c[1]), .O(n13121));
    defparam rd_addr_r_0__bdd_4_lut_11145.LUT_INIT = 16'he4aa;
    SB_DFF i4469_4470 (.Q(\REG.mem_46_5 ), .C(FIFO_CLK_c), .D(n5694));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4466_4467 (.Q(\REG.mem_46_4 ), .C(FIFO_CLK_c), .D(n5693));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4463_4464 (.Q(\REG.mem_46_3 ), .C(FIFO_CLK_c), .D(n5692));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4460_4461 (.Q(\REG.mem_46_2 ), .C(FIFO_CLK_c), .D(n5691));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4457_4458 (.Q(\REG.mem_46_1 ), .C(FIFO_CLK_c), .D(n5690));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4454_4455 (.Q(\REG.mem_46_0 ), .C(FIFO_CLK_c), .D(n5689));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4403_4404 (.Q(\REG.mem_45_15 ), .C(FIFO_CLK_c), .D(n5688));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4400_4401 (.Q(\REG.mem_45_14 ), .C(FIFO_CLK_c), .D(n5687));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4397_4398 (.Q(\REG.mem_45_13 ), .C(FIFO_CLK_c), .D(n5686));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4394_4395 (.Q(\REG.mem_45_12 ), .C(FIFO_CLK_c), .D(n5685));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4391_4392 (.Q(\REG.mem_45_11 ), .C(FIFO_CLK_c), .D(n5684));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4388_4389 (.Q(\REG.mem_45_10 ), .C(FIFO_CLK_c), .D(n5683));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4385_4386 (.Q(\REG.mem_45_9 ), .C(FIFO_CLK_c), .D(n5682));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4382_4383 (.Q(\REG.mem_45_8 ), .C(FIFO_CLK_c), .D(n5681));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4379_4380 (.Q(\REG.mem_45_7 ), .C(FIFO_CLK_c), .D(n5680));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4376_4377 (.Q(\REG.mem_45_6 ), .C(FIFO_CLK_c), .D(n5679));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut (.I0(rd_addr_r_c[1]), .I1(n11861), .I2(n11862), 
            .I3(rd_addr_r_c[2]), .O(n13835));
    defparam rd_addr_r_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n13121_bdd_4_lut (.I0(n13121), .I1(\REG.mem_53_3 ), .I2(\REG.mem_52_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11119));
    defparam n13121_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13835_bdd_4_lut (.I0(n13835), .I1(n11859), .I2(n11858), .I3(rd_addr_r_c[2]), 
            .O(n11025));
    defparam n13835_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4373_4374 (.Q(\REG.mem_45_5 ), .C(FIFO_CLK_c), .D(n5678));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11745 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_6 ), 
            .I2(\REG.mem_39_6 ), .I3(rd_addr_r_c[1]), .O(n13829));
    defparam rd_addr_r_0__bdd_4_lut_11745.LUT_INIT = 16'he4aa;
    SB_LUT4 i3984_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_27_5 ), .O(n5367));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3984_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3983_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_27_4 ), .O(n5366));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3983_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10742 (.I0(rd_addr_r_c[1]), .I1(n11897), 
            .I2(n11898), .I3(rd_addr_r_c[2]), .O(n12467));
    defparam rd_addr_r_1__bdd_4_lut_10742.LUT_INIT = 16'he4aa;
    SB_LUT4 n13829_bdd_4_lut (.I0(n13829), .I1(\REG.mem_37_6 ), .I2(\REG.mem_36_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11407));
    defparam n13829_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12467_bdd_4_lut (.I0(n12467), .I1(n11886), .I2(n11885), .I3(rd_addr_r_c[2]), 
            .O(n12470));
    defparam n12467_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4370_4371 (.Q(\REG.mem_45_4 ), .C(FIFO_CLK_c), .D(n5677));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11140 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_11 ), 
            .I2(\REG.mem_31_11 ), .I3(rd_addr_r_c[1]), .O(n13115));
    defparam rd_addr_r_0__bdd_4_lut_11140.LUT_INIT = 16'he4aa;
    SB_DFF i4367_4368 (.Q(\REG.mem_45_3 ), .C(FIFO_CLK_c), .D(n5676));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13115_bdd_4_lut (.I0(n13115), .I1(\REG.mem_29_11 ), .I2(\REG.mem_28_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11668));
    defparam n13115_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10607 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_5 ), 
            .I2(\REG.mem_43_5 ), .I3(rd_addr_r_c[1]), .O(n12461));
    defparam rd_addr_r_0__bdd_4_lut_10607.LUT_INIT = 16'he4aa;
    SB_DFF i4364_4365 (.Q(\REG.mem_45_2 ), .C(FIFO_CLK_c), .D(n5675));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4361_4362 (.Q(\REG.mem_45_1 ), .C(FIFO_CLK_c), .D(n5674));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4358_4359 (.Q(\REG.mem_45_0 ), .C(FIFO_CLK_c), .D(n5673));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wr_grey_sync_r__i6 (.Q(wr_grey_sync_r[6]), .C(FIFO_CLK_c), .D(n5672));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFF i4307_4308 (.Q(\REG.mem_44_15 ), .C(FIFO_CLK_c), .D(n5671));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4304_4305 (.Q(\REG.mem_44_14 ), .C(FIFO_CLK_c), .D(n5670));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4301_4302 (.Q(\REG.mem_44_13 ), .C(FIFO_CLK_c), .D(n5669));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4298_4299 (.Q(\REG.mem_44_12 ), .C(FIFO_CLK_c), .D(n5668));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4295_4296 (.Q(\REG.mem_44_11 ), .C(FIFO_CLK_c), .D(n5666));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4292_4293 (.Q(\REG.mem_44_10 ), .C(FIFO_CLK_c), .D(n5665));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4289_4290 (.Q(\REG.mem_44_9 ), .C(FIFO_CLK_c), .D(n5664));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4286_4287 (.Q(\REG.mem_44_8 ), .C(FIFO_CLK_c), .D(n5662));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4283_4284 (.Q(\REG.mem_44_7 ), .C(FIFO_CLK_c), .D(n5661));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_4__bdd_4_lut (.I0(rd_addr_r_c[4]), .I1(n11392), .I2(n11401), 
            .I3(rd_addr_r_c[5]), .O(n13823));
    defparam rd_addr_r_4__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11135 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_1 ), 
            .I2(\REG.mem_55_1 ), .I3(rd_addr_r_c[1]), .O(n13109));
    defparam rd_addr_r_0__bdd_4_lut_11135.LUT_INIT = 16'he4aa;
    SB_LUT4 i3982_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_27_3 ), .O(n5365));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3982_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13109_bdd_4_lut (.I0(n13109), .I1(\REG.mem_53_1 ), .I2(\REG.mem_52_1 ), 
            .I3(rd_addr_r_c[1]), .O(n13112));
    defparam n13109_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3981_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_27_2 ), .O(n5364));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3981_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3980_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_27_1 ), .O(n5363));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3980_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i4280_4281 (.Q(\REG.mem_44_6 ), .C(FIFO_CLK_c), .D(n5660));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4277_4278 (.Q(\REG.mem_44_5 ), .C(FIFO_CLK_c), .D(n5659));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4274_4275 (.Q(\REG.mem_44_4 ), .C(FIFO_CLK_c), .D(n5658));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4271_4272 (.Q(\REG.mem_44_3 ), .C(FIFO_CLK_c), .D(n5657));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4268_4269 (.Q(\REG.mem_44_2 ), .C(FIFO_CLK_c), .D(n5656));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4265_4266 (.Q(\REG.mem_44_1 ), .C(FIFO_CLK_c), .D(n5655));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4262_4263 (.Q(\REG.mem_44_0 ), .C(FIFO_CLK_c), .D(n5654));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4211_4212 (.Q(\REG.mem_43_15 ), .C(FIFO_CLK_c), .D(n5653));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4208_4209 (.Q(\REG.mem_43_14 ), .C(FIFO_CLK_c), .D(n5652));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4205_4206 (.Q(\REG.mem_43_13 ), .C(FIFO_CLK_c), .D(n5651));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4202_4203 (.Q(\REG.mem_43_12 ), .C(FIFO_CLK_c), .D(n5650));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4199_4200 (.Q(\REG.mem_43_11 ), .C(FIFO_CLK_c), .D(n5649));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4196_4197 (.Q(\REG.mem_43_10 ), .C(FIFO_CLK_c), .D(n5648));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4193_4194 (.Q(\REG.mem_43_9 ), .C(FIFO_CLK_c), .D(n5647));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4190_4191 (.Q(\REG.mem_43_8 ), .C(FIFO_CLK_c), .D(n5646));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4187_4188 (.Q(\REG.mem_43_7 ), .C(FIFO_CLK_c), .D(n5645));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4184_4185 (.Q(\REG.mem_43_6 ), .C(FIFO_CLK_c), .D(n5644));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3979_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_27_0 ), .O(n5362));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3979_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12461_bdd_4_lut (.I0(n12461), .I1(\REG.mem_41_5 ), .I2(\REG.mem_40_5 ), 
            .I3(rd_addr_r_c[1]), .O(n12464));
    defparam n12461_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13823_bdd_4_lut (.I0(n13823), .I1(n11383), .I2(n12320), .I3(rd_addr_r_c[5]), 
            .O(\REG.out_raw_31__N_559 [9]));
    defparam n13823_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_6 (.CI(n10093), .I0(wp_sync_w[4]), 
            .I1(n1[4]), .CO(n10094));
    SB_LUT4 i4010_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_28_15 ), .O(n5393));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4010_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4009_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_28_14 ), .O(n5392));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4009_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4008_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_28_13 ), .O(n5391));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4008_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_5_lut (.I0(GND_net), .I1(wp_sync_w[3]), 
            .I2(n1[3]), .I3(n10092), .O(rd_sig_diff0_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11730 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_1 ), 
            .I2(\REG.mem_23_1 ), .I3(rd_addr_r_c[1]), .O(n13817));
    defparam rd_addr_r_0__bdd_4_lut_11730.LUT_INIT = 16'he4aa;
    SB_LUT4 i4007_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_28_12 ), .O(n5390));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4007_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_6__I_0_151_2_lut (.I0(GND_net), .I1(rd_addr_r[0]), 
            .I2(GND_net), .I3(VCC_net), .O(\rd_addr_p1_w[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_5 (.CI(n10092), .I0(wp_sync_w[3]), 
            .I1(n1[3]), .CO(n10093));
    SB_LUT4 n13817_bdd_4_lut (.I0(n13817), .I1(\REG.mem_21_1 ), .I2(\REG.mem_20_1 ), 
            .I3(rd_addr_r_c[1]), .O(n11419));
    defparam n13817_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11130 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_11 ), 
            .I2(\REG.mem_35_11 ), .I3(rd_addr_r_c[1]), .O(n13103));
    defparam rd_addr_r_0__bdd_4_lut_11130.LUT_INIT = 16'he4aa;
    SB_DFF i4181_4182 (.Q(\REG.mem_43_5 ), .C(FIFO_CLK_c), .D(n5643));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13103_bdd_4_lut (.I0(n13103), .I1(\REG.mem_33_11 ), .I2(\REG.mem_32_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11674));
    defparam n13103_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4178_4179 (.Q(\REG.mem_43_4 ), .C(FIFO_CLK_c), .D(n5642));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4175_4176 (.Q(\REG.mem_43_3 ), .C(FIFO_CLK_c), .D(n5641));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4172_4173 (.Q(\REG.mem_43_2 ), .C(FIFO_CLK_c), .D(n5640));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4169_4170 (.Q(\REG.mem_43_1 ), .C(FIFO_CLK_c), .D(n5639));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4166_4167 (.Q(\REG.mem_43_0 ), .C(FIFO_CLK_c), .D(n5638));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4115_4116 (.Q(\REG.mem_42_15 ), .C(FIFO_CLK_c), .D(n5637));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4112_4113 (.Q(\REG.mem_42_14 ), .C(FIFO_CLK_c), .D(n5636));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4109_4110 (.Q(\REG.mem_42_13 ), .C(FIFO_CLK_c), .D(n5635));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4106_4107 (.Q(\REG.mem_42_12 ), .C(FIFO_CLK_c), .D(n5634));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4103_4104 (.Q(\REG.mem_42_11 ), .C(FIFO_CLK_c), .D(n5633));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4100_4101 (.Q(\REG.mem_42_10 ), .C(FIFO_CLK_c), .D(n5632));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4097_4098 (.Q(\REG.mem_42_9 ), .C(FIFO_CLK_c), .D(n5631));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4094_4095 (.Q(\REG.mem_42_8 ), .C(FIFO_CLK_c), .D(n5630));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4091_4092 (.Q(\REG.mem_42_7 ), .C(FIFO_CLK_c), .D(n5629));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF \genblk16.rd_prev_r_132  (.Q(\genblk16.rd_prev_r ), .C(SLM_CLK_c), 
           .D(n4916));   // src/fifo_dc_32_lut_gen.v(751[29] 761[32])
    SB_LUT4 i4006_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_28_11 ), .O(n5389));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4006_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10539 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_15 ), 
            .I2(\REG.mem_43_15 ), .I3(rd_addr_r_c[1]), .O(n12389));
    defparam rd_addr_r_0__bdd_4_lut_10539.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10642 (.I0(rd_addr_r_c[2]), .I1(n11302), 
            .I2(n12434), .I3(rd_addr_r_c[3]), .O(n12455));
    defparam rd_addr_r_2__bdd_4_lut_10642.LUT_INIT = 16'he4aa;
    SB_LUT4 n12455_bdd_4_lut (.I0(n12455), .I1(n11230), .I2(n12416), .I3(rd_addr_r_c[3]), 
            .O(n12458));
    defparam n12455_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10592 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_6 ), 
            .I2(\REG.mem_31_6 ), .I3(rd_addr_r_c[1]), .O(n12449));
    defparam rd_addr_r_0__bdd_4_lut_10592.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11720 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_2 ), 
            .I2(\REG.mem_23_2 ), .I3(rd_addr_r_c[1]), .O(n13811));
    defparam rd_addr_r_0__bdd_4_lut_11720.LUT_INIT = 16'he4aa;
    SB_LUT4 n12449_bdd_4_lut (.I0(n12449), .I1(\REG.mem_29_6 ), .I2(\REG.mem_28_6 ), 
            .I3(rd_addr_r_c[1]), .O(n12452));
    defparam n12449_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11125 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_11 ), 
            .I2(\REG.mem_39_11 ), .I3(rd_addr_r_c[1]), .O(n13097));
    defparam rd_addr_r_0__bdd_4_lut_11125.LUT_INIT = 16'he4aa;
    SB_LUT4 n13097_bdd_4_lut (.I0(n13097), .I1(\REG.mem_37_11 ), .I2(\REG.mem_36_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11677));
    defparam n13097_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i167_168 (.Q(\REG.mem_1_11 ), .C(FIFO_CLK_c), .D(n4915));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i152_153 (.Q(\REG.mem_1_6 ), .C(FIFO_CLK_c), .D(n4914));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4088_4089 (.Q(\REG.mem_42_6 ), .C(FIFO_CLK_c), .D(n5628));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4085_4086 (.Q(\REG.mem_42_5 ), .C(FIFO_CLK_c), .D(n5627));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4082_4083 (.Q(\REG.mem_42_4 ), .C(FIFO_CLK_c), .D(n5626));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4079_4080 (.Q(\REG.mem_42_3 ), .C(FIFO_CLK_c), .D(n5625));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4076_4077 (.Q(\REG.mem_42_2 ), .C(FIFO_CLK_c), .D(n5624));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4073_4074 (.Q(\REG.mem_42_1 ), .C(FIFO_CLK_c), .D(n5623));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4070_4071 (.Q(\REG.mem_42_0 ), .C(FIFO_CLK_c), .D(n5622));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4019_4020 (.Q(\REG.mem_41_15 ), .C(FIFO_CLK_c), .D(n5621));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4016_4017 (.Q(\REG.mem_41_14 ), .C(FIFO_CLK_c), .D(n5620));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4013_4014 (.Q(\REG.mem_41_13 ), .C(FIFO_CLK_c), .D(n5619));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4010_4011 (.Q(\REG.mem_41_12 ), .C(FIFO_CLK_c), .D(n5618));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4007_4008 (.Q(\REG.mem_41_11 ), .C(FIFO_CLK_c), .D(n5617));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4004_4005 (.Q(\REG.mem_41_10 ), .C(FIFO_CLK_c), .D(n5616));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4001_4002 (.Q(\REG.mem_41_9 ), .C(FIFO_CLK_c), .D(n5615));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3998_3999 (.Q(\REG.mem_41_8 ), .C(FIFO_CLK_c), .D(n5614));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3995_3996 (.Q(\REG.mem_41_7 ), .C(FIFO_CLK_c), .D(n5613));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4005_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_28_10 ), .O(n5388));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4005_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4004_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_28_9 ), .O(n5387));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4004_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13811_bdd_4_lut (.I0(n13811), .I1(\REG.mem_21_2 ), .I2(\REG.mem_20_2 ), 
            .I3(rd_addr_r_c[1]), .O(n13814));
    defparam n13811_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11510 (.I0(rd_addr_r_c[2]), .I1(n12830), 
            .I2(n12770), .I3(rd_addr_r_c[3]), .O(n13091));
    defparam rd_addr_r_2__bdd_4_lut_11510.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10582 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_2 ), 
            .I2(\REG.mem_3_2 ), .I3(rd_addr_r_c[1]), .O(n12443));
    defparam rd_addr_r_0__bdd_4_lut_10582.LUT_INIT = 16'he4aa;
    SB_LUT4 n12443_bdd_4_lut (.I0(n12443), .I1(\REG.mem_1_2 ), .I2(\REG.mem_0_2 ), 
            .I3(rd_addr_r_c[1]), .O(n12446));
    defparam n12443_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i170_171 (.Q(\REG.mem_1_12 ), .C(FIFO_CLK_c), .D(n4912));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3992_3993 (.Q(\REG.mem_41_6 ), .C(FIFO_CLK_c), .D(n5612));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3989_3990 (.Q(\REG.mem_41_5 ), .C(FIFO_CLK_c), .D(n5611));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3986_3987 (.Q(\REG.mem_41_4 ), .C(FIFO_CLK_c), .D(n5610));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3983_3984 (.Q(\REG.mem_41_3 ), .C(FIFO_CLK_c), .D(n5609));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3980_3981 (.Q(\REG.mem_41_2 ), .C(FIFO_CLK_c), .D(n5608));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3977_3978 (.Q(\REG.mem_41_1 ), .C(FIFO_CLK_c), .D(n5607));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3974_3975 (.Q(\REG.mem_41_0 ), .C(FIFO_CLK_c), .D(n5606));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3923_3924 (.Q(\REG.mem_40_15 ), .C(FIFO_CLK_c), .D(n5605));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3920_3921 (.Q(\REG.mem_40_14 ), .C(FIFO_CLK_c), .D(n5604));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3917_3918 (.Q(\REG.mem_40_13 ), .C(FIFO_CLK_c), .D(n5603));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3914_3915 (.Q(\REG.mem_40_12 ), .C(FIFO_CLK_c), .D(n5602));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3911_3912 (.Q(\REG.mem_40_11 ), .C(FIFO_CLK_c), .D(n5601));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3908_3909 (.Q(\REG.mem_40_10 ), .C(FIFO_CLK_c), .D(n5600));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3905_3906 (.Q(\REG.mem_40_9 ), .C(FIFO_CLK_c), .D(n5599));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3902_3903 (.Q(\REG.mem_40_8 ), .C(FIFO_CLK_c), .D(n5598));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3899_3900 (.Q(\REG.mem_40_7 ), .C(FIFO_CLK_c), .D(n5597));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9393_3_lut (.I0(\REG.mem_24_9 ), .I1(\REG.mem_25_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11231));
    defparam i9393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13091_bdd_4_lut (.I0(n13091), .I1(n12854), .I2(n12914), .I3(rd_addr_r_c[3]), 
            .O(n13094));
    defparam n13091_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11715 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_14 ), 
            .I2(\REG.mem_63_14 ), .I3(rd_addr_r_c[1]), .O(n13805));
    defparam rd_addr_r_0__bdd_4_lut_11715.LUT_INIT = 16'he4aa;
    SB_LUT4 i4003_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_28_8 ), .O(n5386));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4003_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY rd_addr_r_6__I_0_151_2 (.CI(VCC_net), .I0(rd_addr_r[0]), .I1(GND_net), 
            .CO(n10139));
    SB_DFF i155_156 (.Q(\REG.mem_1_7 ), .C(FIFO_CLK_c), .D(n4905));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9394_3_lut (.I0(\REG.mem_26_9 ), .I1(\REG.mem_27_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11232));
    defparam i9394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13805_bdd_4_lut (.I0(n13805), .I1(\REG.mem_61_14 ), .I2(\REG.mem_60_14 ), 
            .I3(rd_addr_r_c[1]), .O(n10996));
    defparam n13805_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF wp_sync2_r__i0 (.Q(wp_sync2_r[0]), .C(SLM_CLK_c), .D(n4904));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_LUT4 i4002_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_28_7 ), .O(n5385));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4002_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF wp_sync1_r__i0 (.Q(wp_sync1_r[0]), .C(SLM_CLK_c), .D(n4903));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF i173_174 (.Q(\REG.mem_1_13 ), .C(FIFO_CLK_c), .D(n4902));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rd_addr_r__i0 (.Q(rd_addr_r[0]), .C(SLM_CLK_c), .D(n4901));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF i158_159 (.Q(\REG.mem_1_8 ), .C(FIFO_CLK_c), .D(n4900));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync2_r__i0 (.Q(rp_sync2_r[0]), .C(FIFO_CLK_c), .D(n4899));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF i3896_3897 (.Q(\REG.mem_40_6 ), .C(FIFO_CLK_c), .D(n5596));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11170 (.I0(rd_addr_r_c[3]), .I1(n11567), 
            .I2(n11568), .I3(rd_addr_r_c[4]), .O(n13085));
    defparam rd_addr_r_3__bdd_4_lut_11170.LUT_INIT = 16'he4aa;
    SB_DFF i3893_3894 (.Q(\REG.mem_40_5 ), .C(FIFO_CLK_c), .D(n5595));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3890_3891 (.Q(\REG.mem_40_4 ), .C(FIFO_CLK_c), .D(n5594));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3887_3888 (.Q(\REG.mem_40_3 ), .C(FIFO_CLK_c), .D(n5593));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3884_3885 (.Q(\REG.mem_40_2 ), .C(FIFO_CLK_c), .D(n5592));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3881_3882 (.Q(\REG.mem_40_1 ), .C(FIFO_CLK_c), .D(n5591));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3878_3879 (.Q(\REG.mem_40_0 ), .C(FIFO_CLK_c), .D(n5590));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3827_3828 (.Q(\REG.mem_39_15 ), .C(FIFO_CLK_c), .D(n5589));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3824_3825 (.Q(\REG.mem_39_14 ), .C(FIFO_CLK_c), .D(n5588));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3821_3822 (.Q(\REG.mem_39_13 ), .C(FIFO_CLK_c), .D(n5587));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3818_3819 (.Q(\REG.mem_39_12 ), .C(FIFO_CLK_c), .D(n5586));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3815_3816 (.Q(\REG.mem_39_11 ), .C(FIFO_CLK_c), .D(n5585));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3812_3813 (.Q(\REG.mem_39_10 ), .C(FIFO_CLK_c), .D(n5584));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3809_3810 (.Q(\REG.mem_39_9 ), .C(FIFO_CLK_c), .D(n5583));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3806_3807 (.Q(\REG.mem_39_8 ), .C(FIFO_CLK_c), .D(n5582));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3803_3804 (.Q(\REG.mem_39_7 ), .C(FIFO_CLK_c), .D(n5581));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync1_r__i0 (.Q(rp_sync1_r[0]), .C(FIFO_CLK_c), .D(n4898));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_LUT4 rd_addr_r_3__bdd_4_lut (.I0(rd_addr_r_c[3]), .I1(n12680), .I2(n11022), 
            .I3(rd_addr_r_c[4]), .O(n13799));
    defparam rd_addr_r_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n13799_bdd_4_lut (.I0(n13799), .I1(n11019), .I2(n12674), .I3(rd_addr_r_c[4]), 
            .O(n13802));
    defparam n13799_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut (.I0(wr_sig_diff0_w[0]), .I1(wr_sig_diff0_w[1]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_23));   // src/fifo_dc_32_lut_gen.v(403[38:87])
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10577 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_1 ), 
            .I2(\REG.mem_15_1 ), .I3(rd_addr_r_c[1]), .O(n12431));
    defparam rd_addr_r_0__bdd_4_lut_10577.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut (.I0(DEBUG_5_c), .I1(wr_sig_diff0_w[3]), .I2(n6_adj_23), 
            .I3(wr_sig_diff0_w[2]), .O(n2_adj_22));   // src/fifo_dc_32_lut_gen.v(403[38:87])
    defparam i1_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 n12431_bdd_4_lut (.I0(n12431), .I1(\REG.mem_13_1 ), .I2(\REG.mem_12_1 ), 
            .I3(rd_addr_r_c[1]), .O(n12434));
    defparam n12431_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13085_bdd_4_lut (.I0(n13085), .I1(n11553), .I2(n13040), .I3(rd_addr_r_c[4]), 
            .O(n13088));
    defparam n13085_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11710 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_3 ), 
            .I2(\REG.mem_3_3 ), .I3(rd_addr_r_c[1]), .O(n13793));
    defparam rd_addr_r_0__bdd_4_lut_11710.LUT_INIT = 16'he4aa;
    SB_LUT4 n13793_bdd_4_lut (.I0(n13793), .I1(\REG.mem_1_3 ), .I2(\REG.mem_0_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11035));
    defparam n13793_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut (.I0(wr_sig_diff0_w[2]), .I1(wr_sig_diff0_w[1]), .I2(wr_sig_diff0_w[0]), 
            .I3(GND_net), .O(n10254));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9114_4_lut (.I0(dc32_fifo_almost_full), .I1(n10925), .I2(n10254), 
            .I3(wr_sig_diff0_w[3]), .O(n10951));
    defparam i9114_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11110 (.I0(rd_addr_r_c[3]), .I1(n13046), 
            .I2(n11559), .I3(rd_addr_r_c[4]), .O(n13079));
    defparam rd_addr_r_3__bdd_4_lut_11110.LUT_INIT = 16'he4aa;
    SB_LUT4 n13079_bdd_4_lut (.I0(n13079), .I1(n11550), .I2(n13034), .I3(rd_addr_r_c[4]), 
            .O(n13082));
    defparam n13079_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4001_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_28_6 ), .O(n5384));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4001_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3800_3801 (.Q(\REG.mem_39_6 ), .C(FIFO_CLK_c), .D(n5580));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3797_3798 (.Q(\REG.mem_39_5 ), .C(FIFO_CLK_c), .D(n5579));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4000_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_28_5 ), .O(n5383));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4000_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3794_3795 (.Q(\REG.mem_39_4 ), .C(FIFO_CLK_c), .D(n5578));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3791_3792 (.Q(\REG.mem_39_3 ), .C(FIFO_CLK_c), .D(n5577));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3788_3789 (.Q(\REG.mem_39_2 ), .C(FIFO_CLK_c), .D(n5576));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3785_3786 (.Q(\REG.mem_39_1 ), .C(FIFO_CLK_c), .D(n5575));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3782_3783 (.Q(\REG.mem_39_0 ), .C(FIFO_CLK_c), .D(n5573));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3731_3732 (.Q(\REG.mem_38_15 ), .C(FIFO_CLK_c), .D(n5572));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3728_3729 (.Q(\REG.mem_38_14 ), .C(FIFO_CLK_c), .D(n5571));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3725_3726 (.Q(\REG.mem_38_13 ), .C(FIFO_CLK_c), .D(n5570));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3722_3723 (.Q(\REG.mem_38_12 ), .C(FIFO_CLK_c), .D(n5569));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3719_3720 (.Q(\REG.mem_38_11 ), .C(FIFO_CLK_c), .D(n5568));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3716_3717 (.Q(\REG.mem_38_10 ), .C(FIFO_CLK_c), .D(n5567));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3713_3714 (.Q(\REG.mem_38_9 ), .C(FIFO_CLK_c), .D(n5566));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3710_3711 (.Q(\REG.mem_38_8 ), .C(FIFO_CLK_c), .D(n5565));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3707_3708 (.Q(\REG.mem_38_7 ), .C(FIFO_CLK_c), .D(n5564));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3999_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_28_4 ), .O(n5382));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3999_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3998_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_28_3 ), .O(n5381));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3998_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3997_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_28_2 ), .O(n5380));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3997_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3996_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_28_1 ), .O(n5379));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3996_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3995_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_28_0 ), .O(n5378));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3995_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4026_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_29_15 ), .O(n5409));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4026_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4025_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_29_14 ), .O(n5408));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4025_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12389_bdd_4_lut (.I0(n12389), .I1(\REG.mem_41_15 ), .I2(\REG.mem_40_15 ), 
            .I3(rd_addr_r_c[1]), .O(n12392));
    defparam n12389_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4024_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_29_13 ), .O(n5407));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4024_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4023_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_29_12 ), .O(n5406));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4023_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4022_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_29_11 ), .O(n5405));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4022_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4021_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_29_10 ), .O(n5404));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4021_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10499 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_5 ), 
            .I2(\REG.mem_47_5 ), .I3(rd_addr_r_c[1]), .O(n12341));
    defparam rd_addr_r_0__bdd_4_lut_10499.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11700 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_13 ), 
            .I2(\REG.mem_43_13 ), .I3(rd_addr_r_c[1]), .O(n13787));
    defparam rd_addr_r_0__bdd_4_lut_11700.LUT_INIT = 16'he4aa;
    SB_LUT4 n13787_bdd_4_lut (.I0(n13787), .I1(\REG.mem_41_13 ), .I2(\REG.mem_40_13 ), 
            .I3(rd_addr_r_c[1]), .O(n11440));
    defparam n13787_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4020_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_29_9 ), .O(n5403));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4020_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3704_3705 (.Q(\REG.mem_38_6 ), .C(FIFO_CLK_c), .D(n5563));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3701_3702 (.Q(\REG.mem_38_5 ), .C(FIFO_CLK_c), .D(n5562));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3698_3699 (.Q(\REG.mem_38_4 ), .C(FIFO_CLK_c), .D(n5561));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3695_3696 (.Q(\REG.mem_38_3 ), .C(FIFO_CLK_c), .D(n5560));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3692_3693 (.Q(\REG.mem_38_2 ), .C(FIFO_CLK_c), .D(n5559));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3689_3690 (.Q(\REG.mem_38_1 ), .C(FIFO_CLK_c), .D(n5558));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3686_3687 (.Q(\REG.mem_38_0 ), .C(FIFO_CLK_c), .D(n5556));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3635_3636 (.Q(\REG.mem_37_15 ), .C(FIFO_CLK_c), .D(n5555));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3632_3633 (.Q(\REG.mem_37_14 ), .C(FIFO_CLK_c), .D(n5554));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3629_3630 (.Q(\REG.mem_37_13 ), .C(FIFO_CLK_c), .D(n5553));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3626_3627 (.Q(\REG.mem_37_12 ), .C(FIFO_CLK_c), .D(n5552));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3623_3624 (.Q(\REG.mem_37_11 ), .C(FIFO_CLK_c), .D(n5551));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3620_3621 (.Q(\REG.mem_37_10 ), .C(FIFO_CLK_c), .D(n5550));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3617_3618 (.Q(\REG.mem_37_9 ), .C(FIFO_CLK_c), .D(n5549));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11155 (.I0(rd_addr_r_c[1]), .I1(n11504), 
            .I2(n11505), .I3(rd_addr_r_c[2]), .O(n13073));
    defparam rd_addr_r_1__bdd_4_lut_11155.LUT_INIT = 16'he4aa;
    SB_LUT4 n13073_bdd_4_lut (.I0(n13073), .I1(n11475), .I2(n11474), .I3(rd_addr_r_c[2]), 
            .O(n13076));
    defparam n13073_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11695 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_13 ), 
            .I2(\REG.mem_27_13 ), .I3(rd_addr_r_c[1]), .O(n13781));
    defparam rd_addr_r_0__bdd_4_lut_11695.LUT_INIT = 16'he4aa;
    SB_LUT4 i4019_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_29_8 ), .O(n5402));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4019_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13781_bdd_4_lut (.I0(n13781), .I1(\REG.mem_25_13 ), .I2(\REG.mem_24_13 ), 
            .I3(rd_addr_r_c[1]), .O(n13784));
    defparam n13781_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4018_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_29_7 ), .O(n5401));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4018_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \REG.out_raw__i16  (.Q(\REG.out_raw[15] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [15]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i15  (.Q(\REG.out_raw[14] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [14]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i14  (.Q(\REG.out_raw[13] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [13]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i13  (.Q(\REG.out_raw[12] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [12]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i12  (.Q(\REG.out_raw[11] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [11]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFF i3614_3615 (.Q(\REG.mem_37_8 ), .C(FIFO_CLK_c), .D(n5548));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3611_3612 (.Q(\REG.mem_37_7 ), .C(FIFO_CLK_c), .D(n5547));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3608_3609 (.Q(\REG.mem_37_6 ), .C(FIFO_CLK_c), .D(n5546));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3605_3606 (.Q(\REG.mem_37_5 ), .C(FIFO_CLK_c), .D(n5545));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3602_3603 (.Q(\REG.mem_37_4 ), .C(FIFO_CLK_c), .D(n5544));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3599_3600 (.Q(\REG.mem_37_3 ), .C(FIFO_CLK_c), .D(n5543));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3596_3597 (.Q(\REG.mem_37_2 ), .C(FIFO_CLK_c), .D(n5542));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3593_3594 (.Q(\REG.mem_37_1 ), .C(FIFO_CLK_c), .D(n5541));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3590_3591 (.Q(\REG.mem_37_0 ), .C(FIFO_CLK_c), .D(n5540));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11100 (.I0(rd_addr_r_c[1]), .I1(n11519), 
            .I2(n11520), .I3(rd_addr_r_c[2]), .O(n13067));
    defparam rd_addr_r_1__bdd_4_lut_11100.LUT_INIT = 16'he4aa;
    SB_LUT4 i4017_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_29_6 ), .O(n5400));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4017_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \REG.out_raw__i11  (.Q(\REG.out_raw[10] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [10]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i10  (.Q(\REG.out_raw[9] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [9]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i9  (.Q(\REG.out_raw[8] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [8]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFSR wr_grey_sync_r__i5 (.Q(wr_grey_sync_r[5]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[5]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFE \REG.out_raw__i8  (.Q(\REG.out_raw[7] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [7]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFSR wr_grey_sync_r__i4 (.Q(wr_grey_sync_r[4]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[4]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFE \REG.out_raw__i7  (.Q(\REG.out_raw[6] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [6]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFSR wr_grey_sync_r__i3 (.Q(wr_grey_sync_r[3]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[3]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFE \REG.out_raw__i6  (.Q(\REG.out_raw[5] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [5]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFSR wr_grey_sync_r__i2 (.Q(wr_grey_sync_r[2]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[2]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFE \REG.out_raw__i5  (.Q(\REG.out_raw[4] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [4]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFSR wr_grey_sync_r__i1 (.Q(wr_grey_sync_r[1]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[1]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFE \REG.out_raw__i4  (.Q(\REG.out_raw[3] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [3]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i3  (.Q(\REG.out_raw[2] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [2]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i2  (.Q(\REG.out_raw[1] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [1]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11690 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_2 ), 
            .I2(\REG.mem_43_2 ), .I3(rd_addr_r_c[1]), .O(n13775));
    defparam rd_addr_r_0__bdd_4_lut_11690.LUT_INIT = 16'he4aa;
    SB_LUT4 i4016_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_29_5 ), .O(n5399));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4016_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3539_3540 (.Q(\REG.mem_36_15 ), .C(FIFO_CLK_c), .D(n5526));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3536_3537 (.Q(\REG.mem_36_14 ), .C(FIFO_CLK_c), .D(n5525));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3533_3534 (.Q(\REG.mem_36_13 ), .C(FIFO_CLK_c), .D(n5524));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3530_3531 (.Q(\REG.mem_36_12 ), .C(FIFO_CLK_c), .D(n5523));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3527_3528 (.Q(\REG.mem_36_11 ), .C(FIFO_CLK_c), .D(n5522));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3524_3525 (.Q(\REG.mem_36_10 ), .C(FIFO_CLK_c), .D(n5521));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3521_3522 (.Q(\REG.mem_36_9 ), .C(FIFO_CLK_c), .D(n5520));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3518_3519 (.Q(\REG.mem_36_8 ), .C(FIFO_CLK_c), .D(n5519));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3515_3516 (.Q(\REG.mem_36_7 ), .C(FIFO_CLK_c), .D(n5518));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3512_3513 (.Q(\REG.mem_36_6 ), .C(FIFO_CLK_c), .D(n5517));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3509_3510 (.Q(\REG.mem_36_5 ), .C(FIFO_CLK_c), .D(n5516));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4015_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_29_4 ), .O(n5398));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4015_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10017_3_lut (.I0(\REG.mem_48_8 ), .I1(\REG.mem_49_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11855));
    defparam i10017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_141_8_lut (.I0(GND_net), .I1(wr_grey_sync_r[6]), 
            .I2(GND_net), .I3(n10138), .O(wr_addr_p1_w[6])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_4_lut (.I0(GND_net), .I1(wp_sync_w[2]), 
            .I2(n1[2]), .I3(n10091), .O(\rd_sig_diff0_w[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4014_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_29_3 ), .O(n5397));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4014_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3506_3507 (.Q(\REG.mem_36_4 ), .C(FIFO_CLK_c), .D(n5515));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3503_3504 (.Q(\REG.mem_36_3 ), .C(FIFO_CLK_c), .D(n5514));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3500_3501 (.Q(\REG.mem_36_2 ), .C(FIFO_CLK_c), .D(n5513));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3497_3498 (.Q(\REG.mem_36_1 ), .C(FIFO_CLK_c), .D(n5512));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3494_3495 (.Q(\REG.mem_36_0 ), .C(FIFO_CLK_c), .D(n5511));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3443_3444 (.Q(\REG.mem_35_15 ), .C(FIFO_CLK_c), .D(n5507));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4013_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_29_2 ), .O(n5396));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4013_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3440_3441 (.Q(\REG.mem_35_14 ), .C(FIFO_CLK_c), .D(n5506));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3437_3438 (.Q(\REG.mem_35_13 ), .C(FIFO_CLK_c), .D(n5505));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3434_3435 (.Q(\REG.mem_35_12 ), .C(FIFO_CLK_c), .D(n5504));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3431_3432 (.Q(\REG.mem_35_11 ), .C(FIFO_CLK_c), .D(n5503));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3428_3429 (.Q(\REG.mem_35_10 ), .C(FIFO_CLK_c), .D(n5502));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3425_3426 (.Q(\REG.mem_35_9 ), .C(FIFO_CLK_c), .D(n5501));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3422_3423 (.Q(\REG.mem_35_8 ), .C(FIFO_CLK_c), .D(n5500));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10018_3_lut (.I0(\REG.mem_50_8 ), .I1(\REG.mem_51_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11856));
    defparam i10018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13775_bdd_4_lut (.I0(n13775), .I1(\REG.mem_41_2 ), .I2(\REG.mem_40_2 ), 
            .I3(rd_addr_r_c[1]), .O(n13778));
    defparam n13775_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_4 (.CI(n10091), .I0(wp_sync_w[2]), 
            .I1(n1[2]), .CO(n10092));
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_3_lut (.I0(GND_net), .I1(wp_sync_w[1]), 
            .I2(n1[1]), .I3(n10090), .O(\rd_sig_diff0_w[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10027_3_lut (.I0(\REG.mem_54_8 ), .I1(\REG.mem_55_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11865));
    defparam i10027_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i3419_3420 (.Q(\REG.mem_35_7 ), .C(FIFO_CLK_c), .D(n5499));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3416_3417 (.Q(\REG.mem_35_6 ), .C(FIFO_CLK_c), .D(n5498));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3413_3414 (.Q(\REG.mem_35_5 ), .C(FIFO_CLK_c), .D(n5497));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3410_3411 (.Q(\REG.mem_35_4 ), .C(FIFO_CLK_c), .D(n5496));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3407_3408 (.Q(\REG.mem_35_3 ), .C(FIFO_CLK_c), .D(n5495));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3404_3405 (.Q(\REG.mem_35_2 ), .C(FIFO_CLK_c), .D(n5494));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3401_3402 (.Q(\REG.mem_35_1 ), .C(FIFO_CLK_c), .D(n5493));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3398_3399 (.Q(\REG.mem_35_0 ), .C(FIFO_CLK_c), .D(n5492));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3347_3348 (.Q(\REG.mem_34_15 ), .C(FIFO_CLK_c), .D(n5490));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3344_3345 (.Q(\REG.mem_34_14 ), .C(FIFO_CLK_c), .D(n5489));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3341_3342 (.Q(\REG.mem_34_13 ), .C(FIFO_CLK_c), .D(n5488));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3338_3339 (.Q(\REG.mem_34_12 ), .C(FIFO_CLK_c), .D(n5487));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3335_3336 (.Q(\REG.mem_34_11 ), .C(FIFO_CLK_c), .D(n5486));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3332_3333 (.Q(\REG.mem_34_10 ), .C(FIFO_CLK_c), .D(n5485));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3329_3330 (.Q(\REG.mem_34_9 ), .C(FIFO_CLK_c), .D(n5484));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4012_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_29_1 ), .O(n5395));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4012_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4011_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_29_0 ), .O(n5394));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4011_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4042_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_30_15 ), .O(n5425));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4042_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10026_3_lut (.I0(\REG.mem_52_8 ), .I1(\REG.mem_53_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11864));
    defparam i10026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4041_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_30_14 ), .O(n5424));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4041_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4040_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_30_13 ), .O(n5423));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4040_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4039_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_30_12 ), .O(n5422));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4039_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4038_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_30_11 ), .O(n5421));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4038_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11735 (.I0(rd_addr_r_c[1]), .I1(n11441), 
            .I2(n11442), .I3(rd_addr_r_c[2]), .O(n13769));
    defparam rd_addr_r_1__bdd_4_lut_11735.LUT_INIT = 16'he4aa;
    SB_LUT4 n13067_bdd_4_lut (.I0(n13067), .I1(n11517), .I2(n11516), .I3(rd_addr_r_c[2]), 
            .O(n13070));
    defparam n13067_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i3326_3327 (.Q(\REG.mem_34_8 ), .C(FIFO_CLK_c), .D(n5483));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3323_3324 (.Q(\REG.mem_34_7 ), .C(FIFO_CLK_c), .D(n5482));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3320_3321 (.Q(\REG.mem_34_6 ), .C(FIFO_CLK_c), .D(n5481));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3317_3318 (.Q(\REG.mem_34_5 ), .C(FIFO_CLK_c), .D(n5480));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3314_3315 (.Q(\REG.mem_34_4 ), .C(FIFO_CLK_c), .D(n5479));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3311_3312 (.Q(\REG.mem_34_3 ), .C(FIFO_CLK_c), .D(n5478));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3308_3309 (.Q(\REG.mem_34_2 ), .C(FIFO_CLK_c), .D(n5477));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3305_3306 (.Q(\REG.mem_34_1 ), .C(FIFO_CLK_c), .D(n5476));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3302_3303 (.Q(\REG.mem_34_0 ), .C(FIFO_CLK_c), .D(n5474));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3251_3252 (.Q(\REG.mem_33_15 ), .C(FIFO_CLK_c), .D(n5473));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3248_3249 (.Q(\REG.mem_33_14 ), .C(FIFO_CLK_c), .D(n5472));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3245_3246 (.Q(\REG.mem_33_13 ), .C(FIFO_CLK_c), .D(n5471));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3242_3243 (.Q(\REG.mem_33_12 ), .C(FIFO_CLK_c), .D(n5470));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3239_3240 (.Q(\REG.mem_33_11 ), .C(FIFO_CLK_c), .D(n5469));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3236_3237 (.Q(\REG.mem_33_10 ), .C(FIFO_CLK_c), .D(n5468));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4037_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_30_10 ), .O(n5420));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4037_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13769_bdd_4_lut (.I0(n13769), .I1(n11394), .I2(n11393), .I3(rd_addr_r_c[2]), 
            .O(n12020));
    defparam n13769_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4036_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_30_9 ), .O(n5419));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4036_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11095 (.I0(rd_addr_r_c[1]), .I1(n11429), 
            .I2(n11430), .I3(rd_addr_r_c[2]), .O(n13061));
    defparam rd_addr_r_1__bdd_4_lut_11095.LUT_INIT = 16'he4aa;
    SB_LUT4 i4035_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_30_8 ), .O(n5418));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4035_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11685 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_3 ), 
            .I2(\REG.mem_7_3 ), .I3(rd_addr_r_c[1]), .O(n13763));
    defparam rd_addr_r_0__bdd_4_lut_11685.LUT_INIT = 16'he4aa;
    SB_LUT4 n13763_bdd_4_lut (.I0(n13763), .I1(\REG.mem_5_3 ), .I2(\REG.mem_4_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11041));
    defparam n13763_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i3233_3234 (.Q(\REG.mem_33_9 ), .C(FIFO_CLK_c), .D(n5467));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3230_3231 (.Q(\REG.mem_33_8 ), .C(FIFO_CLK_c), .D(n5466));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3227_3228 (.Q(\REG.mem_33_7 ), .C(FIFO_CLK_c), .D(n5465));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3224_3225 (.Q(\REG.mem_33_6 ), .C(FIFO_CLK_c), .D(n5464));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3221_3222 (.Q(\REG.mem_33_5 ), .C(FIFO_CLK_c), .D(n5463));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3218_3219 (.Q(\REG.mem_33_4 ), .C(FIFO_CLK_c), .D(n5462));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3215_3216 (.Q(\REG.mem_33_3 ), .C(FIFO_CLK_c), .D(n5461));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3212_3213 (.Q(\REG.mem_33_2 ), .C(FIFO_CLK_c), .D(n5460));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3209_3210 (.Q(\REG.mem_33_1 ), .C(FIFO_CLK_c), .D(n5459));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3206_3207 (.Q(\REG.mem_33_0 ), .C(FIFO_CLK_c), .D(n5458));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3155_3156 (.Q(\REG.mem_32_15 ), .C(FIFO_CLK_c), .D(n5457));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3152_3153 (.Q(\REG.mem_32_14 ), .C(FIFO_CLK_c), .D(n5456));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3149_3150 (.Q(\REG.mem_32_13 ), .C(FIFO_CLK_c), .D(n5455));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3146_3147 (.Q(\REG.mem_32_12 ), .C(FIFO_CLK_c), .D(n5454));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3143_3144 (.Q(\REG.mem_32_11 ), .C(FIFO_CLK_c), .D(n5453));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13061_bdd_4_lut (.I0(n13061), .I1(n11412), .I2(n11411), .I3(rd_addr_r_c[2]), 
            .O(n13064));
    defparam n13061_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4034_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_30_7 ), .O(n5417));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4034_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11090 (.I0(rd_addr_r_c[1]), .I1(n11285), 
            .I2(n11286), .I3(rd_addr_r_c[2]), .O(n13055));
    defparam rd_addr_r_1__bdd_4_lut_11090.LUT_INIT = 16'he4aa;
    SB_DFF i3140_3141 (.Q(\REG.mem_32_10 ), .C(FIFO_CLK_c), .D(n5452));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4033_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_30_6 ), .O(n5416));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4033_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3137_3138 (.Q(\REG.mem_32_9 ), .C(FIFO_CLK_c), .D(n5451));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3134_3135 (.Q(\REG.mem_32_8 ), .C(FIFO_CLK_c), .D(n5450));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3131_3132 (.Q(\REG.mem_32_7 ), .C(FIFO_CLK_c), .D(n5449));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3128_3129 (.Q(\REG.mem_32_6 ), .C(FIFO_CLK_c), .D(n5448));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3125_3126 (.Q(\REG.mem_32_5 ), .C(FIFO_CLK_c), .D(n5447));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3122_3123 (.Q(\REG.mem_32_4 ), .C(FIFO_CLK_c), .D(n5446));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3119_3120 (.Q(\REG.mem_32_3 ), .C(FIFO_CLK_c), .D(n5445));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3116_3117 (.Q(\REG.mem_32_2 ), .C(FIFO_CLK_c), .D(n5444));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3113_3114 (.Q(\REG.mem_32_1 ), .C(FIFO_CLK_c), .D(n5443));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3110_3111 (.Q(\REG.mem_32_0 ), .C(FIFO_CLK_c), .D(n5442));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3059_3060 (.Q(\REG.mem_31_15 ), .C(FIFO_CLK_c), .D(n5441));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3056_3057 (.Q(\REG.mem_31_14 ), .C(FIFO_CLK_c), .D(n5440));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3053_3054 (.Q(\REG.mem_31_13 ), .C(FIFO_CLK_c), .D(n5439));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3050_3051 (.Q(\REG.mem_31_12 ), .C(FIFO_CLK_c), .D(n5438));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3047_3048 (.Q(\REG.mem_31_11 ), .C(FIFO_CLK_c), .D(n5437));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11675 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_1 ), 
            .I2(\REG.mem_27_1 ), .I3(rd_addr_r_c[1]), .O(n13757));
    defparam rd_addr_r_0__bdd_4_lut_11675.LUT_INIT = 16'he4aa;
    SB_LUT4 n13757_bdd_4_lut (.I0(n13757), .I1(\REG.mem_25_1 ), .I2(\REG.mem_24_1 ), 
            .I3(rd_addr_r_c[1]), .O(n11455));
    defparam n13757_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13055_bdd_4_lut (.I0(n13055), .I1(n11283), .I2(n11282), .I3(rd_addr_r_c[2]), 
            .O(n13058));
    defparam n13055_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i3044_3045 (.Q(\REG.mem_31_10 ), .C(FIFO_CLK_c), .D(n5436));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4032_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_30_5 ), .O(n5415));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4032_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4031_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_30_4 ), .O(n5414));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4031_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i84_2_lut_3_lut (.I0(n36), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n58));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i84_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11085 (.I0(rd_addr_r_c[1]), .I1(n11489), 
            .I2(n11490), .I3(rd_addr_r_c[2]), .O(n13049));
    defparam rd_addr_r_1__bdd_4_lut_11085.LUT_INIT = 16'he4aa;
    SB_LUT4 i4030_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_30_3 ), .O(n5413));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4030_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3041_3042 (.Q(\REG.mem_31_9 ), .C(FIFO_CLK_c), .D(n5435));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3038_3039 (.Q(\REG.mem_31_8 ), .C(FIFO_CLK_c), .D(n5434));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3035_3036 (.Q(\REG.mem_31_7 ), .C(FIFO_CLK_c), .D(n5433));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3032_3033 (.Q(\REG.mem_31_6 ), .C(FIFO_CLK_c), .D(n5432));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3029_3030 (.Q(\REG.mem_31_5 ), .C(FIFO_CLK_c), .D(n5431));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3026_3027 (.Q(\REG.mem_31_4 ), .C(FIFO_CLK_c), .D(n5430));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3023_3024 (.Q(\REG.mem_31_3 ), .C(FIFO_CLK_c), .D(n5429));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3020_3021 (.Q(\REG.mem_31_2 ), .C(FIFO_CLK_c), .D(n5428));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3017_3018 (.Q(\REG.mem_31_1 ), .C(FIFO_CLK_c), .D(n5427));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3014_3015 (.Q(\REG.mem_31_0 ), .C(FIFO_CLK_c), .D(n5426));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2963_2964 (.Q(\REG.mem_30_15 ), .C(FIFO_CLK_c), .D(n5425));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2960_2961 (.Q(\REG.mem_30_14 ), .C(FIFO_CLK_c), .D(n5424));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2957_2958 (.Q(\REG.mem_30_13 ), .C(FIFO_CLK_c), .D(n5423));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2954_2955 (.Q(\REG.mem_30_12 ), .C(FIFO_CLK_c), .D(n5422));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2951_2952 (.Q(\REG.mem_30_11 ), .C(FIFO_CLK_c), .D(n5421));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2948_2949 (.Q(\REG.mem_30_10 ), .C(FIFO_CLK_c), .D(n5420));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10044_3_lut (.I0(\REG.mem_48_15 ), .I1(\REG.mem_49_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11882));
    defparam i10044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10045_3_lut (.I0(\REG.mem_50_15 ), .I1(\REG.mem_51_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11883));
    defparam i10045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10057_3_lut (.I0(\REG.mem_54_15 ), .I1(\REG.mem_55_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11895));
    defparam i10057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_inv_0_i7_1_lut (.I0(rp_sync2_r[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_45[6]));   // src/fifo_dc_32_lut_gen.v(212[47:78])
    defparam wr_addr_r_6__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4029_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_30_2 ), .O(n5412));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4029_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13049_bdd_4_lut (.I0(n13049), .I1(n11478), .I2(n11477), .I3(rd_addr_r_c[2]), 
            .O(n13052));
    defparam n13049_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10056_3_lut (.I0(\REG.mem_52_15 ), .I1(\REG.mem_53_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11894));
    defparam i10056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4028_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_30_1 ), .O(n5411));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4028_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11670 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_2 ), 
            .I2(\REG.mem_47_2 ), .I3(rd_addr_r_c[1]), .O(n13751));
    defparam rd_addr_r_0__bdd_4_lut_11670.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11080 (.I0(rd_addr_r_c[1]), .I1(n11450), 
            .I2(n11451), .I3(rd_addr_r_c[2]), .O(n13043));
    defparam rd_addr_r_1__bdd_4_lut_11080.LUT_INIT = 16'he4aa;
    SB_DFF i2945_2946 (.Q(\REG.mem_30_9 ), .C(FIFO_CLK_c), .D(n5419));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2942_2943 (.Q(\REG.mem_30_8 ), .C(FIFO_CLK_c), .D(n5418));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2939_2940 (.Q(\REG.mem_30_7 ), .C(FIFO_CLK_c), .D(n5417));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2936_2937 (.Q(\REG.mem_30_6 ), .C(FIFO_CLK_c), .D(n5416));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2933_2934 (.Q(\REG.mem_30_5 ), .C(FIFO_CLK_c), .D(n5415));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2930_2931 (.Q(\REG.mem_30_4 ), .C(FIFO_CLK_c), .D(n5414));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2927_2928 (.Q(\REG.mem_30_3 ), .C(FIFO_CLK_c), .D(n5413));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2924_2925 (.Q(\REG.mem_30_2 ), .C(FIFO_CLK_c), .D(n5412));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2921_2922 (.Q(\REG.mem_30_1 ), .C(FIFO_CLK_c), .D(n5411));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2918_2919 (.Q(\REG.mem_30_0 ), .C(FIFO_CLK_c), .D(n5410));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2867_2868 (.Q(\REG.mem_29_15 ), .C(FIFO_CLK_c), .D(n5409));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2864_2865 (.Q(\REG.mem_29_14 ), .C(FIFO_CLK_c), .D(n5408));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2861_2862 (.Q(\REG.mem_29_13 ), .C(FIFO_CLK_c), .D(n5407));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2858_2859 (.Q(\REG.mem_29_12 ), .C(FIFO_CLK_c), .D(n5406));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2855_2856 (.Q(\REG.mem_29_11 ), .C(FIFO_CLK_c), .D(n5405));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2852_2853 (.Q(\REG.mem_29_10 ), .C(FIFO_CLK_c), .D(n5404));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13043_bdd_4_lut (.I0(n13043), .I1(n11448), .I2(n11447), .I3(rd_addr_r_c[2]), 
            .O(n13046));
    defparam n13043_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4027_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_30_0 ), .O(n5410));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4027_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13751_bdd_4_lut (.I0(n13751), .I1(\REG.mem_45_2 ), .I2(\REG.mem_44_2 ), 
            .I3(rd_addr_r_c[1]), .O(n13754));
    defparam n13751_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4074_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_32_15 ), .O(n5457));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4074_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4073_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_32_14 ), .O(n5456));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4073_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4072_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_32_13 ), .O(n5455));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4072_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11075 (.I0(rd_addr_r_c[1]), .I1(n11243), 
            .I2(n11244), .I3(rd_addr_r_c[2]), .O(n13037));
    defparam rd_addr_r_1__bdd_4_lut_11075.LUT_INIT = 16'he4aa;
    SB_LUT4 i4071_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_32_12 ), .O(n5454));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4071_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4070_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_32_11 ), .O(n5453));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4070_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4069_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_32_10 ), .O(n5452));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4069_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4068_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_32_9 ), .O(n5451));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4068_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11705 (.I0(rd_addr_r_c[3]), .I1(n11921), 
            .I2(n11922), .I3(rd_addr_r_c[4]), .O(n13745));
    defparam rd_addr_r_3__bdd_4_lut_11705.LUT_INIT = 16'he4aa;
    SB_LUT4 n13745_bdd_4_lut (.I0(n13745), .I1(n11901), .I2(n11900), .I3(rd_addr_r_c[4]), 
            .O(n13748));
    defparam n13745_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4067_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_32_8 ), .O(n5450));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4067_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4066_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_32_7 ), .O(n5449));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4066_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4065_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_32_6 ), .O(n5448));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4065_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4064_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_32_5 ), .O(n5447));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4064_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2849_2850 (.Q(\REG.mem_29_9 ), .C(FIFO_CLK_c), .D(n5403));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2846_2847 (.Q(\REG.mem_29_8 ), .C(FIFO_CLK_c), .D(n5402));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2843_2844 (.Q(\REG.mem_29_7 ), .C(FIFO_CLK_c), .D(n5401));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2840_2841 (.Q(\REG.mem_29_6 ), .C(FIFO_CLK_c), .D(n5400));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2837_2838 (.Q(\REG.mem_29_5 ), .C(FIFO_CLK_c), .D(n5399));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2834_2835 (.Q(\REG.mem_29_4 ), .C(FIFO_CLK_c), .D(n5398));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2831_2832 (.Q(\REG.mem_29_3 ), .C(FIFO_CLK_c), .D(n5397));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2828_2829 (.Q(\REG.mem_29_2 ), .C(FIFO_CLK_c), .D(n5396));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2825_2826 (.Q(\REG.mem_29_1 ), .C(FIFO_CLK_c), .D(n5395));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2822_2823 (.Q(\REG.mem_29_0 ), .C(FIFO_CLK_c), .D(n5394));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2771_2772 (.Q(\REG.mem_28_15 ), .C(FIFO_CLK_c), .D(n5393));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2768_2769 (.Q(\REG.mem_28_14 ), .C(FIFO_CLK_c), .D(n5392));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2765_2766 (.Q(\REG.mem_28_13 ), .C(FIFO_CLK_c), .D(n5391));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2762_2763 (.Q(\REG.mem_28_12 ), .C(FIFO_CLK_c), .D(n5390));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2759_2760 (.Q(\REG.mem_28_11 ), .C(FIFO_CLK_c), .D(n5389));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2756_2757 (.Q(\REG.mem_28_10 ), .C(FIFO_CLK_c), .D(n5388));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2753_2754 (.Q(\REG.mem_28_9 ), .C(FIFO_CLK_c), .D(n5387));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13037_bdd_4_lut (.I0(n13037), .I1(n11202), .I2(n11201), .I3(rd_addr_r_c[2]), 
            .O(n13040));
    defparam n13037_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4063_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_32_4 ), .O(n5446));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4063_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4062_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_32_3 ), .O(n5445));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4062_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11665 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_6 ), 
            .I2(\REG.mem_43_6 ), .I3(rd_addr_r_c[1]), .O(n13739));
    defparam rd_addr_r_0__bdd_4_lut_11665.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i83_2_lut_3_lut (.I0(n36), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n26));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i83_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i4061_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_32_2 ), .O(n5444));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4061_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2750_2751 (.Q(\REG.mem_28_8 ), .C(FIFO_CLK_c), .D(n5386));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4060_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_32_1 ), .O(n5443));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4060_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4059_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_32_0 ), .O(n5442));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4059_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13739_bdd_4_lut (.I0(n13739), .I1(\REG.mem_41_6 ), .I2(\REG.mem_40_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11464));
    defparam n13739_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4622_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_62_15 ), .O(n6005));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4622_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11740 (.I0(rd_addr_r_c[2]), .I1(n12938), 
            .I2(n12812), .I3(rd_addr_r_c[3]), .O(n13733));
    defparam rd_addr_r_2__bdd_4_lut_11740.LUT_INIT = 16'he4aa;
    SB_DFF i2747_2748 (.Q(\REG.mem_28_7 ), .C(FIFO_CLK_c), .D(n5385));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2744_2745 (.Q(\REG.mem_28_6 ), .C(FIFO_CLK_c), .D(n5384));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2741_2742 (.Q(\REG.mem_28_5 ), .C(FIFO_CLK_c), .D(n5383));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2738_2739 (.Q(\REG.mem_28_4 ), .C(FIFO_CLK_c), .D(n5382));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2735_2736 (.Q(\REG.mem_28_3 ), .C(FIFO_CLK_c), .D(n5381));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2732_2733 (.Q(\REG.mem_28_2 ), .C(FIFO_CLK_c), .D(n5380));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2729_2730 (.Q(\REG.mem_28_1 ), .C(FIFO_CLK_c), .D(n5379));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2726_2727 (.Q(\REG.mem_28_0 ), .C(FIFO_CLK_c), .D(n5378));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2675_2676 (.Q(\REG.mem_27_15 ), .C(FIFO_CLK_c), .D(n5377));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2672_2673 (.Q(\REG.mem_27_14 ), .C(FIFO_CLK_c), .D(n5376));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2669_2670 (.Q(\REG.mem_27_13 ), .C(FIFO_CLK_c), .D(n5375));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2666_2667 (.Q(\REG.mem_27_12 ), .C(FIFO_CLK_c), .D(n5374));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2663_2664 (.Q(\REG.mem_27_11 ), .C(FIFO_CLK_c), .D(n5373));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2660_2661 (.Q(\REG.mem_27_10 ), .C(FIFO_CLK_c), .D(n5372));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2657_2658 (.Q(\REG.mem_27_9 ), .C(FIFO_CLK_c), .D(n5371));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2654_2655 (.Q(\REG.mem_27_8 ), .C(FIFO_CLK_c), .D(n5370));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i134_135 (.Q(\REG.mem_1_0 ), .C(FIFO_CLK_c), .D(n4884));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11070 (.I0(rd_addr_r_c[1]), .I1(n11423), 
            .I2(n11424), .I3(rd_addr_r_c[2]), .O(n13031));
    defparam rd_addr_r_1__bdd_4_lut_11070.LUT_INIT = 16'he4aa;
    SB_LUT4 i4621_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_62_14 ), .O(n6004));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4621_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13733_bdd_4_lut (.I0(n13733), .I1(n13112), .I2(n13214), .I3(rd_addr_r_c[3]), 
            .O(n11941));
    defparam n13733_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13031_bdd_4_lut (.I0(n13031), .I1(n11415), .I2(n11414), .I3(rd_addr_r_c[2]), 
            .O(n13034));
    defparam n13031_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4620_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_62_13 ), .O(n6003));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4620_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11655 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_0 ), 
            .I2(\REG.mem_47_0 ), .I3(rd_addr_r_c[1]), .O(n13727));
    defparam rd_addr_r_0__bdd_4_lut_11655.LUT_INIT = 16'he4aa;
    SB_DFF i2651_2652 (.Q(\REG.mem_27_7 ), .C(FIFO_CLK_c), .D(n5369));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2648_2649 (.Q(\REG.mem_27_6 ), .C(FIFO_CLK_c), .D(n5368));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2645_2646 (.Q(\REG.mem_27_5 ), .C(FIFO_CLK_c), .D(n5367));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2642_2643 (.Q(\REG.mem_27_4 ), .C(FIFO_CLK_c), .D(n5366));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2639_2640 (.Q(\REG.mem_27_3 ), .C(FIFO_CLK_c), .D(n5365));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2636_2637 (.Q(\REG.mem_27_2 ), .C(FIFO_CLK_c), .D(n5364));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2633_2634 (.Q(\REG.mem_27_1 ), .C(FIFO_CLK_c), .D(n5363));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2630_2631 (.Q(\REG.mem_27_0 ), .C(FIFO_CLK_c), .D(n5362));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2579_2580 (.Q(\REG.mem_26_15 ), .C(FIFO_CLK_c), .D(n5361));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2576_2577 (.Q(\REG.mem_26_14 ), .C(FIFO_CLK_c), .D(n5360));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2573_2574 (.Q(\REG.mem_26_13 ), .C(FIFO_CLK_c), .D(n5359));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2570_2571 (.Q(\REG.mem_26_12 ), .C(FIFO_CLK_c), .D(n5358));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2567_2568 (.Q(\REG.mem_26_11 ), .C(FIFO_CLK_c), .D(n5357));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2564_2565 (.Q(\REG.mem_26_10 ), .C(FIFO_CLK_c), .D(n5356));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2561_2562 (.Q(\REG.mem_26_9 ), .C(FIFO_CLK_c), .D(n5355));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2558_2559 (.Q(\REG.mem_26_8 ), .C(FIFO_CLK_c), .D(n5354));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2555_2556 (.Q(\REG.mem_26_7 ), .C(FIFO_CLK_c), .D(n5353));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4619_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_62_12 ), .O(n6002));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4619_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2552_2553 (.Q(\REG.mem_26_6 ), .C(FIFO_CLK_c), .D(n5352));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4618_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_62_11 ), .O(n6001));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4618_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4617_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_62_10 ), .O(n6000));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4617_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13727_bdd_4_lut (.I0(n13727), .I1(\REG.mem_45_0 ), .I2(\REG.mem_44_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11947));
    defparam n13727_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut (.I0(dc32_fifo_almost_full), .I1(DEBUG_1_c_c), .I2(GND_net), 
            .I3(GND_net), .O(write_to_dc32_fifo_latched_N_425));   // src/fifo_dc_32_lut_gen.v(410[29] 422[32])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11105 (.I0(rd_addr_r_c[3]), .I1(n13010), 
            .I2(n11472), .I3(rd_addr_r_c[4]), .O(n13025));
    defparam rd_addr_r_3__bdd_4_lut_11105.LUT_INIT = 16'he4aa;
    SB_DFF i2549_2550 (.Q(\REG.mem_26_5 ), .C(FIFO_CLK_c), .D(n5351));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4616_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_62_9 ), .O(n5999));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4616_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2546_2547 (.Q(\REG.mem_26_4 ), .C(FIFO_CLK_c), .D(n5350));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2543_2544 (.Q(\REG.mem_26_3 ), .C(FIFO_CLK_c), .D(n5349));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2540_2541 (.Q(\REG.mem_26_2 ), .C(FIFO_CLK_c), .D(n5348));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2537_2538 (.Q(\REG.mem_26_1 ), .C(FIFO_CLK_c), .D(n5347));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2534_2535 (.Q(\REG.mem_26_0 ), .C(FIFO_CLK_c), .D(n5346));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2483_2484 (.Q(\REG.mem_25_15 ), .C(FIFO_CLK_c), .D(n5345));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2480_2481 (.Q(\REG.mem_25_14 ), .C(FIFO_CLK_c), .D(n5344));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2477_2478 (.Q(\REG.mem_25_13 ), .C(FIFO_CLK_c), .D(n5343));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2474_2475 (.Q(\REG.mem_25_12 ), .C(FIFO_CLK_c), .D(n5342));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2471_2472 (.Q(\REG.mem_25_11 ), .C(FIFO_CLK_c), .D(n5341));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2468_2469 (.Q(\REG.mem_25_10 ), .C(FIFO_CLK_c), .D(n5340));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2465_2466 (.Q(\REG.mem_25_9 ), .C(FIFO_CLK_c), .D(n5339));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2462_2463 (.Q(\REG.mem_25_8 ), .C(FIFO_CLK_c), .D(n5338));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2459_2460 (.Q(\REG.mem_25_7 ), .C(FIFO_CLK_c), .D(n5337));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2456_2457 (.Q(\REG.mem_25_6 ), .C(FIFO_CLK_c), .D(n5336));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2453_2454 (.Q(\REG.mem_25_5 ), .C(FIFO_CLK_c), .D(n5335));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12341_bdd_4_lut (.I0(n12341), .I1(\REG.mem_45_5 ), .I2(\REG.mem_44_5 ), 
            .I3(rd_addr_r_c[1]), .O(n12344));
    defparam n12341_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4615_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_62_8 ), .O(n5998));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4615_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4614_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_62_7 ), .O(n5997));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4614_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11645 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_2 ), 
            .I2(\REG.mem_59_2 ), .I3(rd_addr_r_c[1]), .O(n13721));
    defparam rd_addr_r_0__bdd_4_lut_11645.LUT_INIT = 16'he4aa;
    SB_LUT4 n13025_bdd_4_lut (.I0(n13025), .I1(n11460), .I2(n12986), .I3(rd_addr_r_c[4]), 
            .O(n13028));
    defparam n13025_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i1_1_lut (.I0(rd_addr_r[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_DFF i2450_2451 (.Q(\REG.mem_25_4 ), .C(FIFO_CLK_c), .D(n5334));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2447_2448 (.Q(\REG.mem_25_3 ), .C(FIFO_CLK_c), .D(n5333));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i2_1_lut (.I0(rd_addr_r_c[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4613_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_62_6 ), .O(n5996));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4613_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13721_bdd_4_lut (.I0(n13721), .I1(\REG.mem_57_2 ), .I2(\REG.mem_56_2 ), 
            .I3(rd_addr_r_c[1]), .O(n13724));
    defparam n13721_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11065 (.I0(rd_addr_r_c[1]), .I1(n11402), 
            .I2(n11403), .I3(rd_addr_r_c[2]), .O(n13019));
    defparam rd_addr_r_1__bdd_4_lut_11065.LUT_INIT = 16'he4aa;
    SB_LUT4 i4612_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_62_5 ), .O(n5995));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4612_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13019_bdd_4_lut (.I0(n13019), .I1(n11385), .I2(n11384), .I3(rd_addr_r_c[2]), 
            .O(n13022));
    defparam n13019_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i2444_2445 (.Q(\REG.mem_25_2 ), .C(FIFO_CLK_c), .D(n5332));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4611_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_62_4 ), .O(n5994));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4611_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2441_2442 (.Q(\REG.mem_25_1 ), .C(FIFO_CLK_c), .D(n5331));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2438_2439 (.Q(\REG.mem_25_0 ), .C(FIFO_CLK_c), .D(n5330));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10113_3_lut (.I0(n13274), .I1(n13190), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11951));
    defparam i10113_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2387_2388 (.Q(\REG.mem_24_15 ), .C(FIFO_CLK_c), .D(n5329));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2384_2385 (.Q(\REG.mem_24_14 ), .C(FIFO_CLK_c), .D(n5328));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2381_2382 (.Q(\REG.mem_24_13 ), .C(FIFO_CLK_c), .D(n5327));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2378_2379 (.Q(\REG.mem_24_12 ), .C(FIFO_CLK_c), .D(n5326));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2375_2376 (.Q(\REG.mem_24_11 ), .C(FIFO_CLK_c), .D(n5325));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2372_2373 (.Q(\REG.mem_24_10 ), .C(FIFO_CLK_c), .D(n5324));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2369_2370 (.Q(\REG.mem_24_9 ), .C(FIFO_CLK_c), .D(n5323));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2366_2367 (.Q(\REG.mem_24_8 ), .C(FIFO_CLK_c), .D(n5322));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2363_2364 (.Q(\REG.mem_24_7 ), .C(FIFO_CLK_c), .D(n5321));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2360_2361 (.Q(\REG.mem_24_6 ), .C(FIFO_CLK_c), .D(n5320));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2357_2358 (.Q(\REG.mem_24_5 ), .C(FIFO_CLK_c), .D(n5319));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2354_2355 (.Q(\REG.mem_24_4 ), .C(FIFO_CLK_c), .D(n5318));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2351_2352 (.Q(\REG.mem_24_3 ), .C(FIFO_CLK_c), .D(n5317));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2348_2349 (.Q(\REG.mem_24_2 ), .C(FIFO_CLK_c), .D(n5316));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2345_2346 (.Q(\REG.mem_24_1 ), .C(FIFO_CLK_c), .D(n5315));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4610_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_62_3 ), .O(n5993));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4610_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11120 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_15 ), 
            .I2(\REG.mem_15_15 ), .I3(rd_addr_r_c[1]), .O(n13013));
    defparam rd_addr_r_0__bdd_4_lut_11120.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11640 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_13 ), 
            .I2(\REG.mem_7_13 ), .I3(rd_addr_r_c[1]), .O(n13715));
    defparam rd_addr_r_0__bdd_4_lut_11640.LUT_INIT = 16'he4aa;
    SB_LUT4 i4609_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_62_2 ), .O(n5992));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4609_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4608_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_62_1 ), .O(n5991));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4608_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10114_3_lut (.I0(n13136), .I1(n13016), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11952));
    defparam i10114_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2342_2343 (.Q(\REG.mem_24_0 ), .C(FIFO_CLK_c), .D(n5307));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2291_2292 (.Q(\REG.mem_23_15 ), .C(FIFO_CLK_c), .D(n5306));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2288_2289 (.Q(\REG.mem_23_14 ), .C(FIFO_CLK_c), .D(n5305));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2285_2286 (.Q(\REG.mem_23_13 ), .C(FIFO_CLK_c), .D(n5304));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2282_2283 (.Q(\REG.mem_23_12 ), .C(FIFO_CLK_c), .D(n5303));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2279_2280 (.Q(\REG.mem_23_11 ), .C(FIFO_CLK_c), .D(n5302));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2276_2277 (.Q(\REG.mem_23_10 ), .C(FIFO_CLK_c), .D(n5301));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2273_2274 (.Q(\REG.mem_23_9 ), .C(FIFO_CLK_c), .D(n5300));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2270_2271 (.Q(\REG.mem_23_8 ), .C(FIFO_CLK_c), .D(n5299));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2267_2268 (.Q(\REG.mem_23_7 ), .C(FIFO_CLK_c), .D(n5298));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2264_2265 (.Q(\REG.mem_23_6 ), .C(FIFO_CLK_c), .D(n5297));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2261_2262 (.Q(\REG.mem_23_5 ), .C(FIFO_CLK_c), .D(n5296));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2258_2259 (.Q(\REG.mem_23_4 ), .C(FIFO_CLK_c), .D(n5295));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2255_2256 (.Q(\REG.mem_23_3 ), .C(FIFO_CLK_c), .D(n5294));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2252_2253 (.Q(\REG.mem_23_2 ), .C(FIFO_CLK_c), .D(n5293));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2249_2250 (.Q(\REG.mem_23_1 ), .C(FIFO_CLK_c), .D(n5292));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2246_2247 (.Q(\REG.mem_23_0 ), .C(FIFO_CLK_c), .D(n5290));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2195_2196 (.Q(\REG.mem_22_15 ), .C(FIFO_CLK_c), .D(n5289));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2192_2193 (.Q(\REG.mem_22_14 ), .C(FIFO_CLK_c), .D(n5288));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2189_2190 (.Q(\REG.mem_22_13 ), .C(FIFO_CLK_c), .D(n5287));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2186_2187 (.Q(\REG.mem_22_12 ), .C(FIFO_CLK_c), .D(n5286));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2183_2184 (.Q(\REG.mem_22_11 ), .C(FIFO_CLK_c), .D(n5285));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4607_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_62_0 ), .O(n5990));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4607_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFSR rd_grey_sync_r__i5 (.Q(\rd_grey_sync_r[5] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[5]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_LUT4 n13715_bdd_4_lut (.I0(n13715), .I1(\REG.mem_5_13 ), .I2(\REG.mem_4_13 ), 
            .I3(rd_addr_r_c[1]), .O(n11959));
    defparam n13715_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR rd_grey_sync_r__i4 (.Q(\rd_grey_sync_r[4] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[4]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i3 (.Q(\rd_grey_sync_r[3] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[3]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i2 (.Q(\rd_grey_sync_r[2] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[2]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i1 (.Q(\rd_grey_sync_r[1] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[1]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFF i2180_2181 (.Q(\REG.mem_22_10 ), .C(FIFO_CLK_c), .D(n5284));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2177_2178 (.Q(\REG.mem_22_9 ), .C(FIFO_CLK_c), .D(n5283));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2174_2175 (.Q(\REG.mem_22_8 ), .C(FIFO_CLK_c), .D(n5282));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2171_2172 (.Q(\REG.mem_22_7 ), .C(FIFO_CLK_c), .D(n5281));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2168_2169 (.Q(\REG.mem_22_6 ), .C(FIFO_CLK_c), .D(n5280));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2165_2166 (.Q(\REG.mem_22_5 ), .C(FIFO_CLK_c), .D(n5279));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2162_2163 (.Q(\REG.mem_22_4 ), .C(FIFO_CLK_c), .D(n5278));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2159_2160 (.Q(\REG.mem_22_3 ), .C(FIFO_CLK_c), .D(n5277));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2156_2157 (.Q(\REG.mem_22_2 ), .C(FIFO_CLK_c), .D(n5276));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2153_2154 (.Q(\REG.mem_22_1 ), .C(FIFO_CLK_c), .D(n5275));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2150_2151 (.Q(\REG.mem_22_0 ), .C(FIFO_CLK_c), .D(n5274));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2099_2100 (.Q(\REG.mem_21_15 ), .C(FIFO_CLK_c), .D(n5273));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2096_2097 (.Q(\REG.mem_21_14 ), .C(FIFO_CLK_c), .D(n5272));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2093_2094 (.Q(\REG.mem_21_13 ), .C(FIFO_CLK_c), .D(n5271));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2090_2091 (.Q(\REG.mem_21_12 ), .C(FIFO_CLK_c), .D(n5270));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2087_2088 (.Q(\REG.mem_21_11 ), .C(FIFO_CLK_c), .D(n5269));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_4__bdd_4_lut_11725 (.I0(rd_addr_r_c[4]), .I1(n11905), 
            .I2(n11941), .I3(rd_addr_r_c[5]), .O(n13709));
    defparam rd_addr_r_4__bdd_4_lut_11725.LUT_INIT = 16'he4aa;
    SB_LUT4 n13013_bdd_4_lut (.I0(n13013), .I1(\REG.mem_13_15 ), .I2(\REG.mem_12_15 ), 
            .I3(rd_addr_r_c[1]), .O(n13016));
    defparam n13013_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13709_bdd_4_lut (.I0(n13709), .I1(n12290), .I2(n12458), .I3(rd_addr_r_c[5]), 
            .O(\REG.out_raw_31__N_559 [1]));
    defparam n13709_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i98_2_lut_3_lut_4_lut (.I0(n17_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n51));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i98_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_DFF i2084_2085 (.Q(\REG.mem_21_10 ), .C(FIFO_CLK_c), .D(n5268));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2081_2082 (.Q(\REG.mem_21_9 ), .C(FIFO_CLK_c), .D(n5267));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2078_2079 (.Q(\REG.mem_21_8 ), .C(FIFO_CLK_c), .D(n5266));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2075_2076 (.Q(\REG.mem_21_7 ), .C(FIFO_CLK_c), .D(n5265));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2072_2073 (.Q(\REG.mem_21_6 ), .C(FIFO_CLK_c), .D(n5264));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2069_2070 (.Q(\REG.mem_21_5 ), .C(FIFO_CLK_c), .D(n5263));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2066_2067 (.Q(\REG.mem_21_4 ), .C(FIFO_CLK_c), .D(n5262));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2063_2064 (.Q(\REG.mem_21_3 ), .C(FIFO_CLK_c), .D(n5261));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2060_2061 (.Q(\REG.mem_21_2 ), .C(FIFO_CLK_c), .D(n5260));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2057_2058 (.Q(\REG.mem_21_1 ), .C(FIFO_CLK_c), .D(n5259));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2054_2055 (.Q(\REG.mem_21_0 ), .C(FIFO_CLK_c), .D(n5257));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2003_2004 (.Q(\REG.mem_20_15 ), .C(FIFO_CLK_c), .D(n5256));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2000_2001 (.Q(\REG.mem_20_14 ), .C(FIFO_CLK_c), .D(n5255));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1997_1998 (.Q(\REG.mem_20_13 ), .C(FIFO_CLK_c), .D(n5254));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1994_1995 (.Q(\REG.mem_20_12 ), .C(FIFO_CLK_c), .D(n5253));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i97_2_lut_3_lut_4_lut (.I0(n17_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n19));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i97_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i4603_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_61_15 ), .O(n5986));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4603_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4602_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_61_14 ), .O(n5985));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4602_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1991_1992 (.Q(\REG.mem_20_11 ), .C(FIFO_CLK_c), .D(n5252));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11055 (.I0(rd_addr_r_c[1]), .I1(n11204), 
            .I2(n11205), .I3(rd_addr_r_c[2]), .O(n13007));
    defparam rd_addr_r_1__bdd_4_lut_11055.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11635 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_13 ), 
            .I2(\REG.mem_47_13 ), .I3(rd_addr_r_c[1]), .O(n13703));
    defparam rd_addr_r_0__bdd_4_lut_11635.LUT_INIT = 16'he4aa;
    SB_LUT4 n13703_bdd_4_lut (.I0(n13703), .I1(\REG.mem_45_13 ), .I2(\REG.mem_44_13 ), 
            .I3(rd_addr_r_c[1]), .O(n11482));
    defparam n13703_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13007_bdd_4_lut (.I0(n13007), .I1(n11163), .I2(n11162), .I3(rd_addr_r_c[2]), 
            .O(n13010));
    defparam n13007_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11625 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_2 ), 
            .I2(\REG.mem_63_2 ), .I3(rd_addr_r_c[1]), .O(n13697));
    defparam rd_addr_r_0__bdd_4_lut_11625.LUT_INIT = 16'he4aa;
    SB_LUT4 i4601_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_61_13 ), .O(n5984));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4601_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4600_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_61_12 ), .O(n5983));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4600_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13697_bdd_4_lut (.I0(n13697), .I1(\REG.mem_61_2 ), .I2(\REG.mem_60_2 ), 
            .I3(rd_addr_r_c[1]), .O(n13700));
    defparam n13697_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4599_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_61_11 ), .O(n5982));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4599_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4598_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_61_10 ), .O(n5981));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4598_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4597_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_61_9 ), .O(n5980));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4597_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4596_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_61_8 ), .O(n5979));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4596_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1988_1989 (.Q(\REG.mem_20_10 ), .C(FIFO_CLK_c), .D(n5251));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11620 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_6 ), 
            .I2(\REG.mem_47_6 ), .I3(rd_addr_r_c[1]), .O(n13691));
    defparam rd_addr_r_0__bdd_4_lut_11620.LUT_INIT = 16'he4aa;
    SB_DFF i1985_1986 (.Q(\REG.mem_20_9 ), .C(FIFO_CLK_c), .D(n5250));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1982_1983 (.Q(\REG.mem_20_8 ), .C(FIFO_CLK_c), .D(n5249));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1979_1980 (.Q(\REG.mem_20_7 ), .C(FIFO_CLK_c), .D(n5248));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1976_1977 (.Q(\REG.mem_20_6 ), .C(FIFO_CLK_c), .D(n5247));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1973_1974 (.Q(\REG.mem_20_5 ), .C(FIFO_CLK_c), .D(n5246));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1970_1971 (.Q(\REG.mem_20_4 ), .C(FIFO_CLK_c), .D(n5245));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1967_1968 (.Q(\REG.mem_20_3 ), .C(FIFO_CLK_c), .D(n5244));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1964_1965 (.Q(\REG.mem_20_2 ), .C(FIFO_CLK_c), .D(n5243));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1961_1962 (.Q(\REG.mem_20_1 ), .C(FIFO_CLK_c), .D(n5242));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1958_1959 (.Q(\REG.mem_20_0 ), .C(FIFO_CLK_c), .D(n5241));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1907_1908 (.Q(\REG.mem_19_15 ), .C(FIFO_CLK_c), .D(n5240));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1904_1905 (.Q(\REG.mem_19_14 ), .C(FIFO_CLK_c), .D(n5239));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1901_1902 (.Q(\REG.mem_19_13 ), .C(FIFO_CLK_c), .D(n5238));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1898_1899 (.Q(\REG.mem_19_12 ), .C(FIFO_CLK_c), .D(n5237));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4595_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_61_7 ), .O(n5978));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4595_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4594_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_61_6 ), .O(n5977));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4594_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_r_6__I_0_135_i2_3_lut (.I0(wr_addr_r[1]), .I1(wr_addr_p1_w[1]), 
            .I2(wr_sig_mv_w), .I3(GND_net), .O(\wr_addr_nxt_c[1] ));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_6__I_0_135_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11050 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_12 ), 
            .I2(\REG.mem_35_12 ), .I3(rd_addr_r_c[1]), .O(n13001));
    defparam rd_addr_r_0__bdd_4_lut_11050.LUT_INIT = 16'he4aa;
    SB_LUT4 i4593_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_61_5 ), .O(n5976));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4593_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4592_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_61_4 ), .O(n5975));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4592_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13691_bdd_4_lut (.I0(n13691), .I1(\REG.mem_45_6 ), .I2(\REG.mem_44_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11485));
    defparam n13691_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13001_bdd_4_lut (.I0(n13001), .I1(\REG.mem_33_12 ), .I2(\REG.mem_32_12 ), 
            .I3(rd_addr_r_c[1]), .O(n13004));
    defparam n13001_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4591_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_61_3 ), .O(n5974));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4591_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4590_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_61_2 ), .O(n5973));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4590_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4090_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_33_15 ), .O(n5473));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4090_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11040 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_0 ), 
            .I2(\REG.mem_11_0 ), .I3(rd_addr_r_c[1]), .O(n12995));
    defparam rd_addr_r_0__bdd_4_lut_11040.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11615 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_3 ), 
            .I2(\REG.mem_11_3 ), .I3(rd_addr_r_c[1]), .O(n13685));
    defparam rd_addr_r_0__bdd_4_lut_11615.LUT_INIT = 16'he4aa;
    SB_DFF i1895_1896 (.Q(\REG.mem_19_11 ), .C(FIFO_CLK_c), .D(n5236));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4589_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_61_1 ), .O(n5972));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4589_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4588_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_61_0 ), .O(n5971));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4588_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1892_1893 (.Q(\REG.mem_19_10 ), .C(FIFO_CLK_c), .D(n5235));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1889_1890 (.Q(\REG.mem_19_9 ), .C(FIFO_CLK_c), .D(n5234));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1886_1887 (.Q(\REG.mem_19_8 ), .C(FIFO_CLK_c), .D(n5233));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1883_1884 (.Q(\REG.mem_19_7 ), .C(FIFO_CLK_c), .D(n5232));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1880_1881 (.Q(\REG.mem_19_6 ), .C(FIFO_CLK_c), .D(n5231));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1877_1878 (.Q(\REG.mem_19_5 ), .C(FIFO_CLK_c), .D(n5230));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1874_1875 (.Q(\REG.mem_19_4 ), .C(FIFO_CLK_c), .D(n5229));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1871_1872 (.Q(\REG.mem_19_3 ), .C(FIFO_CLK_c), .D(n5228));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1868_1869 (.Q(\REG.mem_19_2 ), .C(FIFO_CLK_c), .D(n5227));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1865_1866 (.Q(\REG.mem_19_1 ), .C(FIFO_CLK_c), .D(n5226));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1862_1863 (.Q(\REG.mem_19_0 ), .C(FIFO_CLK_c), .D(n5225));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1811_1812 (.Q(\REG.mem_18_15 ), .C(FIFO_CLK_c), .D(n5224));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1808_1809 (.Q(\REG.mem_18_14 ), .C(FIFO_CLK_c), .D(n5223));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1805_1806 (.Q(\REG.mem_18_13 ), .C(FIFO_CLK_c), .D(n5222));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1802_1803 (.Q(\REG.mem_18_12 ), .C(FIFO_CLK_c), .D(n5221));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1799_1800 (.Q(\REG.mem_18_11 ), .C(FIFO_CLK_c), .D(n5220));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i1_2_lut_adj_28 (.I0(wp_sync2_r[1]), .I1(wp_sync_w[2]), .I2(GND_net), 
            .I3(GND_net), .O(wp_sync_w[1]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_28.LUT_INIT = 16'h6666;
    SB_LUT4 n13685_bdd_4_lut (.I0(n13685), .I1(\REG.mem_9_3 ), .I2(\REG.mem_8_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11044));
    defparam n13685_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12995_bdd_4_lut (.I0(n12995), .I1(\REG.mem_9_0 ), .I2(\REG.mem_8_0 ), 
            .I3(rd_addr_r_c[1]), .O(n12998));
    defparam n12995_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11610 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_13 ), 
            .I2(\REG.mem_11_13 ), .I3(rd_addr_r_c[1]), .O(n13679));
    defparam rd_addr_r_0__bdd_4_lut_11610.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i96_2_lut_3_lut_4_lut (.I0(n15_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n52));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i96_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 n13679_bdd_4_lut (.I0(n13679), .I1(\REG.mem_9_13 ), .I2(\REG.mem_8_13 ), 
            .I3(rd_addr_r_c[1]), .O(n11965));
    defparam n13679_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i95_2_lut_3_lut_4_lut (.I0(n15_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n20));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i95_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_adj_29 (.I0(wp_sync2_r[3]), .I1(wp_sync_w[4]), .I2(GND_net), 
            .I3(GND_net), .O(wp_sync_w[3]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_29.LUT_INIT = 16'h6666;
    SB_DFF i1796_1797 (.Q(\REG.mem_18_10 ), .C(FIFO_CLK_c), .D(n5219));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i1_2_lut_adj_30 (.I0(wp_sync2_r[6]), .I1(wp_sync2_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n4274));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_30.LUT_INIT = 16'h6666;
    SB_DFF i1793_1794 (.Q(\REG.mem_18_9 ), .C(FIFO_CLK_c), .D(n5218));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1790_1791 (.Q(\REG.mem_18_8 ), .C(FIFO_CLK_c), .D(n5217));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1787_1788 (.Q(\REG.mem_18_7 ), .C(FIFO_CLK_c), .D(n5216));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1784_1785 (.Q(\REG.mem_18_6 ), .C(FIFO_CLK_c), .D(n5215));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1781_1782 (.Q(\REG.mem_18_5 ), .C(FIFO_CLK_c), .D(n5214));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1778_1779 (.Q(\REG.mem_18_4 ), .C(FIFO_CLK_c), .D(n5213));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1775_1776 (.Q(\REG.mem_18_3 ), .C(FIFO_CLK_c), .D(n5212));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1772_1773 (.Q(\REG.mem_18_2 ), .C(FIFO_CLK_c), .D(n5211));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1769_1770 (.Q(\REG.mem_18_1 ), .C(FIFO_CLK_c), .D(n5210));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1766_1767 (.Q(\REG.mem_18_0 ), .C(FIFO_CLK_c), .D(n5209));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1715_1716 (.Q(\REG.mem_17_15 ), .C(FIFO_CLK_c), .D(n5208));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1712_1713 (.Q(\REG.mem_17_14 ), .C(FIFO_CLK_c), .D(n5207));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1709_1710 (.Q(\REG.mem_17_13 ), .C(FIFO_CLK_c), .D(n5206));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1706_1707 (.Q(\REG.mem_17_12 ), .C(FIFO_CLK_c), .D(n5205));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1703_1704 (.Q(\REG.mem_17_11 ), .C(FIFO_CLK_c), .D(n5204));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9053_4_lut (.I0(rd_addr_r[0]), .I1(rd_addr_r_c[4]), .I2(wp_sync_w[0]), 
            .I3(wp_sync_w[4]), .O(n10889));
    defparam i9053_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i9062_4_lut (.I0(rd_addr_r_c[5]), .I1(rd_addr_r_c[3]), .I2(n4274), 
            .I3(wp_sync_w[3]), .O(n10899));
    defparam i9062_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11605 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_0 ), 
            .I2(\REG.mem_51_0 ), .I3(rd_addr_r_c[1]), .O(n13673));
    defparam rd_addr_r_0__bdd_4_lut_11605.LUT_INIT = 16'he4aa;
    SB_LUT4 i3567_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_2_5 ), .O(n4950));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3567_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3566_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_2_4 ), .O(n4949));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3566_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3532_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_1_11 ), .O(n4915));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3532_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1700_1701 (.Q(\REG.mem_17_10 ), .C(FIFO_CLK_c), .D(n5203));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13673_bdd_4_lut (.I0(n13673), .I1(\REG.mem_49_0 ), .I2(\REG.mem_48_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11968));
    defparam n13673_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_31 (.I0(rd_addr_p1_w[4]), .I1(wp_sync_w[4]), .I2(GND_net), 
            .I3(GND_net), .O(n4298));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_31.LUT_INIT = 16'h6666;
    SB_LUT4 i3565_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_2_3 ), .O(n4948));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3565_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3564_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_2_2 ), .O(n4947));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3564_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut (.I0(rd_addr_p1_w[5]), .I1(rd_addr_p1_w[3]), .I2(n4274), 
            .I3(wp_sync_w[3]), .O(n10_c));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i3_4_lut.LUT_INIT = 16'h7bde;
    SB_DFF i1697_1698 (.Q(\REG.mem_17_9 ), .C(FIFO_CLK_c), .D(n5202));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3563_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_2_1 ), .O(n4946));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3563_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11600 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_13 ), 
            .I2(\REG.mem_15_13 ), .I3(rd_addr_r_c[1]), .O(n13667));
    defparam rd_addr_r_0__bdd_4_lut_11600.LUT_INIT = 16'he4aa;
    SB_LUT4 i3562_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_2_0 ), .O(n4945));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3562_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_32 (.I0(wp_sync2_r[6]), .I1(rd_addr_p1_w[1]), .I2(rd_addr_p1_w[6]), 
            .I3(wp_sync_w[1]), .O(n8_adj_25));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i1_4_lut_adj_32.LUT_INIT = 16'h7bde;
    SB_LUT4 i5_4_lut (.I0(\rd_addr_p1_w[0] ), .I1(n10_c), .I2(n4298), 
            .I3(wp_sync_w[0]), .O(n12));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i5_4_lut.LUT_INIT = 16'hfdfe;
    SB_DFF i1694_1695 (.Q(\REG.mem_17_8 ), .C(FIFO_CLK_c), .D(n5201));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9147_3_lut (.I0(n10887), .I1(n10899), .I2(n10889), .I3(GND_net), 
            .O(n10985));
    defparam i9147_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3577_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_2_15 ), .O(n4960));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3577_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13667_bdd_4_lut (.I0(n13667), .I1(\REG.mem_13_13 ), .I2(\REG.mem_12_13 ), 
            .I3(rd_addr_r_c[1]), .O(n11971));
    defparam n13667_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11035 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_9 ), 
            .I2(\REG.mem_43_9 ), .I3(rd_addr_r_c[1]), .O(n12989));
    defparam rd_addr_r_0__bdd_4_lut_11035.LUT_INIT = 16'he4aa;
    SB_LUT4 n12989_bdd_4_lut (.I0(n12989), .I1(\REG.mem_41_9 ), .I2(\REG.mem_40_9 ), 
            .I3(rd_addr_r_c[1]), .O(n12992));
    defparam n12989_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11595 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_4 ), 
            .I2(\REG.mem_7_4 ), .I3(rd_addr_r_c[1]), .O(n13661));
    defparam rd_addr_r_0__bdd_4_lut_11595.LUT_INIT = 16'he4aa;
    SB_LUT4 n13661_bdd_4_lut (.I0(n13661), .I1(\REG.mem_5_4 ), .I2(\REG.mem_4_4 ), 
            .I3(rd_addr_r_c[1]), .O(n13664));
    defparam n13661_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11045 (.I0(rd_addr_r_c[1]), .I1(n11072), 
            .I2(n11073), .I3(rd_addr_r_c[2]), .O(n12983));
    defparam rd_addr_r_1__bdd_4_lut_11045.LUT_INIT = 16'he4aa;
    SB_LUT4 i6_4_lut (.I0(rd_addr_p1_w[2]), .I1(n12), .I2(n8_adj_25), 
            .I3(wp_sync_w[2]), .O(n10258));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i6_4_lut.LUT_INIT = 16'hfdfe;
    SB_LUT4 i3576_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_2_14 ), .O(n4959));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3576_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1691_1692 (.Q(\REG.mem_17_7 ), .C(FIFO_CLK_c), .D(n5200));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1688_1689 (.Q(\REG.mem_17_6 ), .C(FIFO_CLK_c), .D(n5199));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1685_1686 (.Q(\REG.mem_17_5 ), .C(FIFO_CLK_c), .D(n5198));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1682_1683 (.Q(\REG.mem_17_4 ), .C(FIFO_CLK_c), .D(n5197));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1679_1680 (.Q(\REG.mem_17_3 ), .C(FIFO_CLK_c), .D(n5196));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1676_1677 (.Q(\REG.mem_17_2 ), .C(FIFO_CLK_c), .D(n5195));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1673_1674 (.Q(\REG.mem_17_1 ), .C(FIFO_CLK_c), .D(n5194));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 empty_nxt_c_I_7_4_lut (.I0(n10258), .I1(n10985), .I2(DEBUG_3_c), 
            .I3(get_next_word), .O(empty_nxt_c_N_629));   // src/fifo_dc_32_lut_gen.v(555[46:103])
    defparam empty_nxt_c_I_7_4_lut.LUT_INIT = 16'h3530;
    SB_DFF i1670_1671 (.Q(\REG.mem_17_0 ), .C(FIFO_CLK_c), .D(n5193));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1619_1620 (.Q(\REG.mem_16_15 ), .C(FIFO_CLK_c), .D(n5188));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1616_1617 (.Q(\REG.mem_16_14 ), .C(FIFO_CLK_c), .D(n5186));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3575_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_2_13 ), .O(n4958));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3575_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9178_3_lut (.I0(n12740), .I1(n12668), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11016));
    defparam i9178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10173_3_lut (.I0(\REG.mem_0_6 ), .I1(\REG.mem_1_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12011));
    defparam i10173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3574_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_2_12 ), .O(n4957));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3574_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1613_1614 (.Q(\REG.mem_16_13 ), .C(FIFO_CLK_c), .D(n5185));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11590 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_8 ), 
            .I2(\REG.mem_7_8 ), .I3(rd_addr_r_c[1]), .O(n13655));
    defparam rd_addr_r_0__bdd_4_lut_11590.LUT_INIT = 16'he4aa;
    SB_LUT4 i10174_3_lut (.I0(\REG.mem_2_6 ), .I1(\REG.mem_3_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12012));
    defparam i10174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4089_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_33_14 ), .O(n5472));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4089_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1610_1611 (.Q(\REG.mem_16_12 ), .C(FIFO_CLK_c), .D(n5184));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3573_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_2_11 ), .O(n4956));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3573_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13655_bdd_4_lut (.I0(n13655), .I1(\REG.mem_5_8 ), .I2(\REG.mem_4_8 ), 
            .I3(rd_addr_r_c[1]), .O(n13658));
    defparam n13655_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3572_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_2_10 ), .O(n4955));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3572_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10534 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_2 ), 
            .I2(\REG.mem_7_2 ), .I3(rd_addr_r_c[1]), .O(n12383));
    defparam rd_addr_r_0__bdd_4_lut_10534.LUT_INIT = 16'he4aa;
    SB_LUT4 i3571_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_2_9 ), .O(n4954));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3571_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12383_bdd_4_lut (.I0(n12383), .I1(\REG.mem_5_2 ), .I2(\REG.mem_4_2 ), 
            .I3(rd_addr_r_c[1]), .O(n12386));
    defparam n12383_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11680 (.I0(rd_addr_r_c[1]), .I1(n11936), 
            .I2(n11937), .I3(rd_addr_r_c[2]), .O(n13649));
    defparam rd_addr_r_1__bdd_4_lut_11680.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10529 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_9 ), 
            .I2(\REG.mem_63_9 ), .I3(rd_addr_r_c[1]), .O(n12377));
    defparam rd_addr_r_0__bdd_4_lut_10529.LUT_INIT = 16'he4aa;
    SB_LUT4 n12377_bdd_4_lut (.I0(n12377), .I1(\REG.mem_61_9 ), .I2(\REG.mem_60_9 ), 
            .I3(rd_addr_r_c[1]), .O(n12380));
    defparam n12377_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3570_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_2_8 ), .O(n4953));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3570_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3569_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_2_7 ), .O(n4952));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3569_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12983_bdd_4_lut (.I0(n12983), .I1(n11037), .I2(n11036), .I3(rd_addr_r_c[2]), 
            .O(n12986));
    defparam n12983_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13649_bdd_4_lut (.I0(n13649), .I1(n11874), .I2(n11873), .I3(rd_addr_r_c[2]), 
            .O(n11049));
    defparam n13649_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3519_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_1_13 ), .O(n4902));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3519_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3568_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_2_6 ), .O(n4951));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3568_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_6__I_0_i1_3_lut (.I0(rd_addr_r[0]), .I1(\rd_addr_p1_w[0] ), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(rd_addr_nxt_c_6__N_498[0]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_6__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1607_1608 (.Q(\REG.mem_16_11 ), .C(FIFO_CLK_c), .D(n5183));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1604_1605 (.Q(\REG.mem_16_10 ), .C(FIFO_CLK_c), .D(n5182));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1601_1602 (.Q(\REG.mem_16_9 ), .C(FIFO_CLK_c), .D(n5181));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1598_1599 (.Q(\REG.mem_16_8 ), .C(FIFO_CLK_c), .D(n5180));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1595_1596 (.Q(\REG.mem_16_7 ), .C(FIFO_CLK_c), .D(n5179));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1592_1593 (.Q(\REG.mem_16_6 ), .C(FIFO_CLK_c), .D(n5178));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1589_1590 (.Q(\REG.mem_16_5 ), .C(FIFO_CLK_c), .D(n5177));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11585 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_1 ), 
            .I2(\REG.mem_31_1 ), .I3(rd_addr_r_c[1]), .O(n13643));
    defparam rd_addr_r_0__bdd_4_lut_11585.LUT_INIT = 16'he4aa;
    SB_LUT4 n13643_bdd_4_lut (.I0(n13643), .I1(\REG.mem_29_1 ), .I2(\REG.mem_28_1 ), 
            .I3(rd_addr_r_c[1]), .O(n11488));
    defparam n13643_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1586_1587 (.Q(\REG.mem_16_4 ), .C(FIFO_CLK_c), .D(n5176));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i137_138 (.Q(\REG.mem_1_1 ), .C(FIFO_CLK_c), .D(n4879));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4088_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_33_13 ), .O(n5471));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4088_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3529_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_1_12 ), .O(n4912));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3529_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11575 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_13 ), 
            .I2(\REG.mem_51_13 ), .I3(rd_addr_r_c[1]), .O(n13637));
    defparam rd_addr_r_0__bdd_4_lut_11575.LUT_INIT = 16'he4aa;
    SB_LUT4 i10029_3_lut (.I0(\REG.mem_16_14 ), .I1(\REG.mem_17_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11867));
    defparam i10029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10030_3_lut (.I0(\REG.mem_18_14 ), .I1(\REG.mem_19_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11868));
    defparam i10030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9702_3_lut (.I0(\REG.mem_0_12 ), .I1(\REG.mem_1_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11540));
    defparam i9702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13637_bdd_4_lut (.I0(n13637), .I1(\REG.mem_49_13 ), .I2(\REG.mem_48_13 ), 
            .I3(rd_addr_r_c[1]), .O(n11500));
    defparam n13637_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9703_3_lut (.I0(\REG.mem_2_12 ), .I1(\REG.mem_3_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11541));
    defparam i9703_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1583_1584 (.Q(\REG.mem_16_3 ), .C(FIFO_CLK_c), .D(n5175));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1580_1581 (.Q(\REG.mem_16_2 ), .C(FIFO_CLK_c), .D(n5174));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1577_1578 (.Q(\REG.mem_16_1 ), .C(FIFO_CLK_c), .D(n5173));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1574_1575 (.Q(\REG.mem_16_0 ), .C(FIFO_CLK_c), .D(n5172));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1523_1524 (.Q(\REG.mem_15_15 ), .C(FIFO_CLK_c), .D(n5169));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1520_1521 (.Q(\REG.mem_15_14 ), .C(FIFO_CLK_c), .D(n5168));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1517_1518 (.Q(\REG.mem_15_13 ), .C(FIFO_CLK_c), .D(n5167));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i106_2_lut_3_lut_4_lut (.I0(n18_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n47));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i106_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11030 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_11 ), 
            .I2(\REG.mem_43_11 ), .I3(rd_addr_r_c[1]), .O(n12977));
    defparam rd_addr_r_0__bdd_4_lut_11030.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11580 (.I0(rd_addr_r_c[1]), .I1(n11927), 
            .I2(n11928), .I3(rd_addr_r_c[2]), .O(n13631));
    defparam rd_addr_r_1__bdd_4_lut_11580.LUT_INIT = 16'he4aa;
    SB_DFF i1514_1515 (.Q(\REG.mem_15_12 ), .C(FIFO_CLK_c), .D(n5166));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i105_2_lut_3_lut_4_lut (.I0(n18_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n15));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i105_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_DFF i1511_1512 (.Q(\REG.mem_15_11 ), .C(FIFO_CLK_c), .D(n5165));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1508_1509 (.Q(\REG.mem_15_10 ), .C(FIFO_CLK_c), .D(n5164));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1505_1506 (.Q(\REG.mem_15_9 ), .C(FIFO_CLK_c), .D(n5163));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1502_1503 (.Q(\REG.mem_15_8 ), .C(FIFO_CLK_c), .D(n5162));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13631_bdd_4_lut (.I0(n13631), .I1(n11919), .I2(n11918), .I3(rd_addr_r_c[2]), 
            .O(n11052));
    defparam n13631_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1499_1500 (.Q(\REG.mem_15_7 ), .C(FIFO_CLK_c), .D(n5161));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3448_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_1_10 ), .O(n4831));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3448_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12977_bdd_4_lut (.I0(n12977), .I1(\REG.mem_41_11 ), .I2(\REG.mem_40_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11692));
    defparam n12977_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1496_1497 (.Q(\REG.mem_15_6 ), .C(FIFO_CLK_c), .D(n5160));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1493_1494 (.Q(\REG.mem_15_5 ), .C(FIFO_CLK_c), .D(n5159));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1490_1491 (.Q(\REG.mem_15_4 ), .C(FIFO_CLK_c), .D(n5158));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1487_1488 (.Q(\REG.mem_15_3 ), .C(FIFO_CLK_c), .D(n5157));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1484_1485 (.Q(\REG.mem_15_2 ), .C(FIFO_CLK_c), .D(n5156));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1481_1482 (.Q(\REG.mem_15_1 ), .C(FIFO_CLK_c), .D(n5155));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11020 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_12 ), 
            .I2(\REG.mem_39_12 ), .I3(rd_addr_r_c[1]), .O(n12971));
    defparam rd_addr_r_0__bdd_4_lut_11020.LUT_INIT = 16'he4aa;
    SB_DFF i1478_1479 (.Q(\REG.mem_15_0 ), .C(FIFO_CLK_c), .D(n5154));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1427_1428 (.Q(\REG.mem_14_15 ), .C(FIFO_CLK_c), .D(n5153));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1424_1425 (.Q(\REG.mem_14_14 ), .C(FIFO_CLK_c), .D(n5152));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4586_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_60_15 ), .O(n5969));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4586_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4585_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_60_14 ), .O(n5968));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4585_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10186_3_lut (.I0(\REG.mem_6_6 ), .I1(\REG.mem_7_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12024));
    defparam i10186_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1421_1422 (.Q(\REG.mem_14_13 ), .C(FIFO_CLK_c), .D(n5151));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1418_1419 (.Q(\REG.mem_14_12 ), .C(FIFO_CLK_c), .D(n5150));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1415_1416 (.Q(\REG.mem_14_11 ), .C(FIFO_CLK_c), .D(n5149));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1412_1413 (.Q(\REG.mem_14_10 ), .C(FIFO_CLK_c), .D(n5148));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1409_1410 (.Q(\REG.mem_14_9 ), .C(FIFO_CLK_c), .D(n5147));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1406_1407 (.Q(\REG.mem_14_8 ), .C(FIFO_CLK_c), .D(n5146));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1403_1404 (.Q(\REG.mem_14_7 ), .C(FIFO_CLK_c), .D(n5145));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1400_1401 (.Q(\REG.mem_14_6 ), .C(FIFO_CLK_c), .D(n5144));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10185_3_lut (.I0(\REG.mem_4_6 ), .I1(\REG.mem_5_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12023));
    defparam i10185_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1397_1398 (.Q(\REG.mem_14_5 ), .C(FIFO_CLK_c), .D(n5143));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4584_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_60_13 ), .O(n5967));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4584_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1394_1395 (.Q(\REG.mem_14_4 ), .C(FIFO_CLK_c), .D(n5142));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11570 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_9 ), 
            .I2(\REG.mem_15_9 ), .I3(rd_addr_r_c[1]), .O(n13625));
    defparam rd_addr_r_0__bdd_4_lut_11570.LUT_INIT = 16'he4aa;
    SB_DFF i1391_1392 (.Q(\REG.mem_14_3 ), .C(FIFO_CLK_c), .D(n5141));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12971_bdd_4_lut (.I0(n12971), .I1(\REG.mem_37_12 ), .I2(\REG.mem_36_12 ), 
            .I3(rd_addr_r_c[1]), .O(n12974));
    defparam n12971_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1388_1389 (.Q(\REG.mem_14_2 ), .C(FIFO_CLK_c), .D(n5140));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1385_1386 (.Q(\REG.mem_14_1 ), .C(FIFO_CLK_c), .D(n5139));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1382_1383 (.Q(\REG.mem_14_0 ), .C(FIFO_CLK_c), .D(n5138));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1331_1332 (.Q(\REG.mem_13_15 ), .C(FIFO_CLK_c), .D(n5137));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1328_1329 (.Q(\REG.mem_13_14 ), .C(FIFO_CLK_c), .D(n5136));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1325_1326 (.Q(\REG.mem_13_13 ), .C(FIFO_CLK_c), .D(n5135));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1322_1323 (.Q(\REG.mem_13_12 ), .C(FIFO_CLK_c), .D(n5134));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1319_1320 (.Q(\REG.mem_13_11 ), .C(FIFO_CLK_c), .D(n5133));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1316_1317 (.Q(\REG.mem_13_10 ), .C(FIFO_CLK_c), .D(n5132));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13625_bdd_4_lut (.I0(n13625), .I1(\REG.mem_13_9 ), .I2(\REG.mem_12_9 ), 
            .I3(rd_addr_r_c[1]), .O(n11176));
    defparam n13625_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1313_1314 (.Q(\REG.mem_13_9 ), .C(FIFO_CLK_c), .D(n5131));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11560 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_8 ), 
            .I2(\REG.mem_27_8 ), .I3(rd_addr_r_c[1]), .O(n13619));
    defparam rd_addr_r_0__bdd_4_lut_11560.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11015 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_11 ), 
            .I2(\REG.mem_47_11 ), .I3(rd_addr_r_c[1]), .O(n12965));
    defparam rd_addr_r_0__bdd_4_lut_11015.LUT_INIT = 16'he4aa;
    SB_LUT4 n12965_bdd_4_lut (.I0(n12965), .I1(\REG.mem_45_11 ), .I2(\REG.mem_44_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11701));
    defparam n12965_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11025 (.I0(rd_addr_r_c[1]), .I1(n11279), 
            .I2(n11280), .I3(rd_addr_r_c[2]), .O(n12959));
    defparam rd_addr_r_1__bdd_4_lut_11025.LUT_INIT = 16'he4aa;
    SB_LUT4 i3450_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_1_9 ), .O(n4833));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3450_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13619_bdd_4_lut (.I0(n13619), .I1(\REG.mem_25_8 ), .I2(\REG.mem_24_8 ), 
            .I3(rd_addr_r_c[1]), .O(n13622));
    defparam n13619_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4583_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_60_12 ), .O(n5966));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4583_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4582_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_60_11 ), .O(n5965));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4582_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4581_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_60_10 ), .O(n5964));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4581_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3484_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_1_14 ), .O(n4867));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3484_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3522_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_1_7 ), .O(n4905));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3522_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12959_bdd_4_lut (.I0(n12959), .I1(n11253), .I2(n11252), .I3(rd_addr_r_c[2]), 
            .O(n12962));
    defparam n12959_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3531_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_1_6 ), .O(n4914));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3531_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4087_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_33_12 ), .O(n5470));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4087_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1310_1311 (.Q(\REG.mem_13_8 ), .C(FIFO_CLK_c), .D(n5130));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4580_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_60_9 ), .O(n5963));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4580_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4579_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_60_8 ), .O(n5962));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4579_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3449_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_1_15 ), .O(n4832));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3449_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11555 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_0 ), 
            .I2(\REG.mem_55_0 ), .I3(rd_addr_r_c[1]), .O(n13613));
    defparam rd_addr_r_0__bdd_4_lut_11555.LUT_INIT = 16'he4aa;
    SB_LUT4 i4578_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_60_7 ), .O(n5961));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4578_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13613_bdd_4_lut (.I0(n13613), .I1(\REG.mem_53_0 ), .I2(\REG.mem_52_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11977));
    defparam n13613_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4577_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_60_6 ), .O(n5960));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4577_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1307_1308 (.Q(\REG.mem_13_7 ), .C(FIFO_CLK_c), .D(n5129));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1304_1305 (.Q(\REG.mem_13_6 ), .C(FIFO_CLK_c), .D(n5128));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1301_1302 (.Q(\REG.mem_13_5 ), .C(FIFO_CLK_c), .D(n5127));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1298_1299 (.Q(\REG.mem_13_4 ), .C(FIFO_CLK_c), .D(n5126));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4576_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_60_5 ), .O(n5959));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4576_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4575_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_60_4 ), .O(n5958));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4575_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1295_1296 (.Q(\REG.mem_13_3 ), .C(FIFO_CLK_c), .D(n5125));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11005 (.I0(rd_addr_r_c[1]), .I1(n11210), 
            .I2(n11211), .I3(rd_addr_r_c[2]), .O(n12953));
    defparam rd_addr_r_1__bdd_4_lut_11005.LUT_INIT = 16'he4aa;
    SB_LUT4 i4574_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_60_3 ), .O(n5957));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4574_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12953_bdd_4_lut (.I0(n12953), .I1(n11187), .I2(n11186), .I3(rd_addr_r_c[2]), 
            .O(n12956));
    defparam n12953_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1292_1293 (.Q(\REG.mem_13_2 ), .C(FIFO_CLK_c), .D(n5124));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11650 (.I0(rd_addr_r_c[2]), .I1(n13298), 
            .I2(n12482), .I3(rd_addr_r_c[3]), .O(n13607));
    defparam rd_addr_r_2__bdd_4_lut_11650.LUT_INIT = 16'he4aa;
    SB_LUT4 n13607_bdd_4_lut (.I0(n13607), .I1(n11977), .I2(n11968), .I3(rd_addr_r_c[3]), 
            .O(n11983));
    defparam n13607_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1289_1290 (.Q(\REG.mem_13_1 ), .C(FIFO_CLK_c), .D(n5123));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3452_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_1_5 ), .O(n4835));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3452_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3454_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_1_4 ), .O(n4837));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3454_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11550 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_8 ), 
            .I2(\REG.mem_11_8 ), .I3(rd_addr_r_c[1]), .O(n13601));
    defparam rd_addr_r_0__bdd_4_lut_11550.LUT_INIT = 16'he4aa;
    SB_LUT4 i10033_3_lut (.I0(\REG.mem_22_14 ), .I1(\REG.mem_23_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11871));
    defparam i10033_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1286_1287 (.Q(\REG.mem_13_0 ), .C(FIFO_CLK_c), .D(n5122));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1235_1236 (.Q(\REG.mem_12_15 ), .C(FIFO_CLK_c), .D(n5121));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1232_1233 (.Q(\REG.mem_12_14 ), .C(FIFO_CLK_c), .D(n5120));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4573_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_60_2 ), .O(n5956));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4573_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1229_1230 (.Q(\REG.mem_12_13 ), .C(FIFO_CLK_c), .D(n5119));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1226_1227 (.Q(\REG.mem_12_12 ), .C(FIFO_CLK_c), .D(n5118));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3478_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_1_3 ), .O(n4861));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3478_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10524 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_6 ), 
            .I2(\REG.mem_35_6 ), .I3(rd_addr_r_c[1]), .O(n12371));
    defparam rd_addr_r_0__bdd_4_lut_10524.LUT_INIT = 16'he4aa;
    SB_LUT4 i3485_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_1_2 ), .O(n4868));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3485_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11010 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_9 ), 
            .I2(\REG.mem_3_9 ), .I3(rd_addr_r_c[1]), .O(n12947));
    defparam rd_addr_r_0__bdd_4_lut_11010.LUT_INIT = 16'he4aa;
    SB_LUT4 n13601_bdd_4_lut (.I0(n13601), .I1(\REG.mem_9_8 ), .I2(\REG.mem_8_8 ), 
            .I3(rd_addr_r_c[1]), .O(n13604));
    defparam n13601_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1223_1224 (.Q(\REG.mem_12_11 ), .C(FIFO_CLK_c), .D(n5117));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12947_bdd_4_lut (.I0(n12947), .I1(\REG.mem_1_9 ), .I2(\REG.mem_0_9 ), 
            .I3(rd_addr_r_c[1]), .O(n11122));
    defparam n12947_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9162_3_lut (.I0(\REG.mem_8_6 ), .I1(\REG.mem_9_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11000));
    defparam i9162_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1220_1221 (.Q(\REG.mem_12_10 ), .C(FIFO_CLK_c), .D(n5116));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9163_3_lut (.I0(\REG.mem_10_6 ), .I1(\REG.mem_11_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11001));
    defparam i9163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4572_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_60_1 ), .O(n5955));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4572_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11115 (.I0(rd_addr_r_c[2]), .I1(n11272), 
            .I2(n12452), .I3(rd_addr_r_c[3]), .O(n12941));
    defparam rd_addr_r_2__bdd_4_lut_11115.LUT_INIT = 16'he4aa;
    SB_LUT4 i3496_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_1_1 ), .O(n4879));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3496_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4571_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_60_0 ), .O(n5954));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4571_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10032_3_lut (.I0(\REG.mem_20_14 ), .I1(\REG.mem_21_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11870));
    defparam i10032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12941_bdd_4_lut (.I0(n12941), .I1(n11197), .I2(n11110), .I3(rd_addr_r_c[3]), 
            .O(n11704));
    defparam n12941_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3501_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_1_0 ), .O(n4884));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3501_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12287_bdd_4_lut (.I0(n12287), .I1(n11419), .I2(n11389), .I3(rd_addr_r_c[3]), 
            .O(n12290));
    defparam n12287_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i61_2_lut_3_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n61_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i61_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i94_2_lut_3_lut_4_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n53));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i94_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i93_2_lut_3_lut_4_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n21));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i93_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11565 (.I0(rd_addr_r_c[1]), .I1(n11432), 
            .I2(n11433), .I3(rd_addr_r_c[2]), .O(n13595));
    defparam rd_addr_r_1__bdd_4_lut_11565.LUT_INIT = 16'he4aa;
    SB_LUT4 n12371_bdd_4_lut (.I0(n12371), .I1(\REG.mem_33_6 ), .I2(\REG.mem_32_6 ), 
            .I3(rd_addr_r_c[1]), .O(n12374));
    defparam n12371_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i13_2_lut_3_lut_4_lut (.I0(wr_sig_mv_w), .I1(wr_addr_r[0]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[1]), .O(n13));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i13_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i3517_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_1_8 ), .O(n4900));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3517_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10995 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_1 ), 
            .I2(\REG.mem_59_1 ), .I3(rd_addr_r_c[1]), .O(n12935));
    defparam rd_addr_r_0__bdd_4_lut_10995.LUT_INIT = 16'he4aa;
    SB_DFF i1217_1218 (.Q(\REG.mem_12_9 ), .C(FIFO_CLK_c), .D(n5115));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1214_1215 (.Q(\REG.mem_12_8 ), .C(FIFO_CLK_c), .D(n5114));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1211_1212 (.Q(\REG.mem_12_7 ), .C(FIFO_CLK_c), .D(n5113));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i14_2_lut_3_lut_4_lut (.I0(wr_sig_mv_w), .I1(wr_addr_r[0]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[1]), .O(n14));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i14_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 n12935_bdd_4_lut (.I0(n12935), .I1(\REG.mem_57_1 ), .I2(\REG.mem_56_1 ), 
            .I3(rd_addr_r_c[1]), .O(n12938));
    defparam n12935_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4561_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_59_15 ), .O(n5944));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4561_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13595_bdd_4_lut (.I0(n13595), .I1(n11421), .I2(n11420), .I3(rd_addr_r_c[2]), 
            .O(n11514));
    defparam n13595_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4560_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_59_14 ), .O(n5943));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4560_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i2_2_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_w[2]), 
            .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[1] ), .O(wr_grey_w[1]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i2_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11545 (.I0(rd_addr_r_c[2]), .I1(n11440), 
            .I2(n11482), .I3(rd_addr_r_c[3]), .O(n13589));
    defparam rd_addr_r_2__bdd_4_lut_11545.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i3_2_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_w[2]), 
            .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[3] ), .O(wr_grey_w[2]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i3_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_DFF i1208_1209 (.Q(\REG.mem_12_6 ), .C(FIFO_CLK_c), .D(n5112));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4661_2_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_w[2]), 
            .I2(wr_sig_mv_w), .I3(reset_per_frame), .O(n6044));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i4661_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 i4559_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_59_13 ), .O(n5942));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4559_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4086_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_33_11 ), .O(n5469));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4086_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4558_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_59_12 ), .O(n5941));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4558_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4557_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_59_11 ), .O(n5940));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4557_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4556_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_59_10 ), .O(n5939));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4556_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13589_bdd_4_lut (.I0(n13589), .I1(n12398), .I2(n13184), .I3(rd_addr_r_c[3]), 
            .O(n11989));
    defparam n13589_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i100_2_lut_3_lut (.I0(n35), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n50));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i100_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10985 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_11 ), 
            .I2(\REG.mem_51_11 ), .I3(rd_addr_r_c[1]), .O(n12929));
    defparam rd_addr_r_0__bdd_4_lut_10985.LUT_INIT = 16'he4aa;
    SB_DFF i1205_1206 (.Q(\REG.mem_12_5 ), .C(FIFO_CLK_c), .D(n5111));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4555_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_59_9 ), .O(n5938));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4555_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4554_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_59_8 ), .O(n5937));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4554_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i99_2_lut_3_lut (.I0(n35), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n18));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i99_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i9718_3_lut (.I0(\REG.mem_6_12 ), .I1(\REG.mem_7_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11556));
    defparam i9718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4553_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_59_7 ), .O(n5936));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4553_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1202_1203 (.Q(\REG.mem_12_4 ), .C(FIFO_CLK_c), .D(n5110));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1199_1200 (.Q(\REG.mem_12_3 ), .C(FIFO_CLK_c), .D(n5109));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4552_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_59_6 ), .O(n5935));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4552_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4551_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_59_5 ), .O(n5934));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4551_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4550_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_59_4 ), .O(n5933));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4550_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4549_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_59_3 ), .O(n5932));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4549_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1196_1197 (.Q(\REG.mem_12_2 ), .C(FIFO_CLK_c), .D(n5108));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i4_2_lut_4_lut (.I0(wr_addr_r[4]), .I1(wr_addr_p1_w[4]), 
            .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[3] ), .O(wr_grey_w[3]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i4_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 n12929_bdd_4_lut (.I0(n12929), .I1(\REG.mem_49_11 ), .I2(\REG.mem_48_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11710));
    defparam n12929_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9717_3_lut (.I0(\REG.mem_4_12 ), .I1(\REG.mem_5_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11555));
    defparam i9717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4548_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_59_2 ), .O(n5931));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4548_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10519 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_2 ), 
            .I2(\REG.mem_11_2 ), .I3(rd_addr_r_c[1]), .O(n12365));
    defparam rd_addr_r_0__bdd_4_lut_10519.LUT_INIT = 16'he4aa;
    SB_LUT4 i4547_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_59_1 ), .O(n5930));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4547_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i5_2_lut_4_lut (.I0(wr_addr_r[4]), .I1(wr_addr_p1_w[4]), 
            .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[5] ), .O(wr_grey_w[4]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i5_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4546_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_59_0 ), .O(n5929));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4546_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1193_1194 (.Q(\REG.mem_12_1 ), .C(FIFO_CLK_c), .D(n5107));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12365_bdd_4_lut (.I0(n12365), .I1(\REG.mem_9_2 ), .I2(\REG.mem_8_2 ), 
            .I3(rd_addr_r_c[1]), .O(n12368));
    defparam n12365_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i92_2_lut_3_lut_4_lut (.I0(n20_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n54));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i92_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i91_2_lut_3_lut_4_lut (.I0(n20_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n22));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i91_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i4659_2_lut_4_lut (.I0(wr_addr_r[4]), .I1(wr_addr_p1_w[4]), 
            .I2(wr_sig_mv_w), .I3(reset_per_frame), .O(n6042));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i4659_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 i4085_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_33_10 ), .O(n5468));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4085_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10980 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_0 ), 
            .I2(\REG.mem_15_0 ), .I3(rd_addr_r_c[1]), .O(n12923));
    defparam rd_addr_r_0__bdd_4_lut_10980.LUT_INIT = 16'he4aa;
    SB_DFF i1190_1191 (.Q(\REG.mem_12_0 ), .C(FIFO_CLK_c), .D(n5106));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i4_2_lut_4_lut (.I0(rd_addr_r_c[4]), 
            .I1(rd_addr_p1_w[4]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_498[3] ), 
            .O(rd_grey_w[3]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i4_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 n12923_bdd_4_lut (.I0(n12923), .I1(\REG.mem_13_0 ), .I2(\REG.mem_12_0 ), 
            .I3(rd_addr_r_c[1]), .O(n12926));
    defparam n12923_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9256_3_lut (.I0(\REG.mem_14_6 ), .I1(\REG.mem_15_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11094));
    defparam i9256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11660 (.I0(rd_addr_r_c[3]), .I1(n13022), 
            .I2(n11514), .I3(rd_addr_r_c[4]), .O(n13583));
    defparam rd_addr_r_3__bdd_4_lut_11660.LUT_INIT = 16'he4aa;
    SB_LUT4 i9255_3_lut (.I0(\REG.mem_12_6 ), .I1(\REG.mem_13_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11093));
    defparam i9255_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1139_1140 (.Q(\REG.mem_11_15 ), .C(FIFO_CLK_c), .D(n5105));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1136_1137 (.Q(\REG.mem_11_14 ), .C(FIFO_CLK_c), .D(n5104));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1133_1134 (.Q(\REG.mem_11_13 ), .C(FIFO_CLK_c), .D(n5103));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1130_1131 (.Q(\REG.mem_11_12 ), .C(FIFO_CLK_c), .D(n5102));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1127_1128 (.Q(\REG.mem_11_11 ), .C(FIFO_CLK_c), .D(n5101));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1124_1125 (.Q(\REG.mem_11_10 ), .C(FIFO_CLK_c), .D(n5100));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1121_1122 (.Q(\REG.mem_11_9 ), .C(FIFO_CLK_c), .D(n5099));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1118_1119 (.Q(\REG.mem_11_8 ), .C(FIFO_CLK_c), .D(n5098));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i140_141 (.Q(\REG.mem_1_2 ), .C(FIFO_CLK_c), .D(n4868));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i176_177 (.Q(\REG.mem_1_14 ), .C(FIFO_CLK_c), .D(n4867));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wr_addr_r__i0 (.Q(wr_addr_r[0]), .C(FIFO_CLK_c), .D(n4866));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF i143_144 (.Q(\REG.mem_1_3 ), .C(FIFO_CLK_c), .D(n4861));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10975 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_12 ), 
            .I2(\REG.mem_43_12 ), .I3(rd_addr_r_c[1]), .O(n12917));
    defparam rd_addr_r_0__bdd_4_lut_10975.LUT_INIT = 16'he4aa;
    SB_LUT4 n13583_bdd_4_lut (.I0(n13583), .I1(n11493), .I2(n11492), .I3(rd_addr_r_c[4]), 
            .O(n13586));
    defparam n13583_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1115_1116 (.Q(\REG.mem_11_7 ), .C(FIFO_CLK_c), .D(n5097));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11540 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_6 ), 
            .I2(\REG.mem_23_6 ), .I3(rd_addr_r_c[1]), .O(n13577));
    defparam rd_addr_r_0__bdd_4_lut_11540.LUT_INIT = 16'he4aa;
    SB_DFF i1112_1113 (.Q(\REG.mem_11_6 ), .C(FIFO_CLK_c), .D(n5096));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1109_1110 (.Q(\REG.mem_11_5 ), .C(FIFO_CLK_c), .D(n5095));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1106_1107 (.Q(\REG.mem_11_4 ), .C(FIFO_CLK_c), .D(n5094));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1103_1104 (.Q(\REG.mem_11_3 ), .C(FIFO_CLK_c), .D(n5093));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1100_1101 (.Q(\REG.mem_11_2 ), .C(FIFO_CLK_c), .D(n5092));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1097_1098 (.Q(\REG.mem_11_1 ), .C(FIFO_CLK_c), .D(n5091));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1094_1095 (.Q(\REG.mem_11_0 ), .C(FIFO_CLK_c), .D(n5090));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1043_1044 (.Q(\REG.mem_10_15 ), .C(FIFO_CLK_c), .D(n5089));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12917_bdd_4_lut (.I0(n12917), .I1(\REG.mem_41_12 ), .I2(\REG.mem_40_12 ), 
            .I3(rd_addr_r_c[1]), .O(n12920));
    defparam n12917_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1040_1041 (.Q(\REG.mem_10_14 ), .C(FIFO_CLK_c), .D(n5088));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10970 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_0 ), 
            .I2(\REG.mem_19_0 ), .I3(rd_addr_r_c[1]), .O(n12911));
    defparam rd_addr_r_0__bdd_4_lut_10970.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i5_2_lut_4_lut (.I0(rd_addr_r_c[4]), 
            .I1(rd_addr_p1_w[4]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_498[5] ), 
            .O(rd_grey_w[4]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i5_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 n13577_bdd_4_lut (.I0(n13577), .I1(\REG.mem_21_6 ), .I2(\REG.mem_20_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11197));
    defparam n13577_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12911_bdd_4_lut (.I0(n12911), .I1(\REG.mem_17_0 ), .I2(\REG.mem_16_0 ), 
            .I3(rd_addr_r_c[1]), .O(n12914));
    defparam n12911_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1037_1038 (.Q(\REG.mem_10_13 ), .C(FIFO_CLK_c), .D(n5087));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1034_1035 (.Q(\REG.mem_10_12 ), .C(FIFO_CLK_c), .D(n5086));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1031_1032 (.Q(\REG.mem_10_11 ), .C(FIFO_CLK_c), .D(n5085));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1028_1029 (.Q(\REG.mem_10_10 ), .C(FIFO_CLK_c), .D(n5084));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1025_1026 (.Q(\REG.mem_10_9 ), .C(FIFO_CLK_c), .D(n5083));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1022_1023 (.Q(\REG.mem_10_8 ), .C(FIFO_CLK_c), .D(n5082));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1019_1020 (.Q(\REG.mem_10_7 ), .C(FIFO_CLK_c), .D(n5081));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1016_1017 (.Q(\REG.mem_10_6 ), .C(FIFO_CLK_c), .D(n5080));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4539_2_lut_4_lut (.I0(rd_addr_r_c[4]), .I1(rd_addr_p1_w[4]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n5922));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4539_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 rd_addr_r_6__I_0_i6_3_lut (.I0(rd_addr_r_c[5]), .I1(rd_addr_p1_w[5]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_6__N_498[5] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_6__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1013_1014 (.Q(\REG.mem_10_5 ), .C(FIFO_CLK_c), .D(n5079));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10965 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_1 ), 
            .I2(\REG.mem_11_1 ), .I3(rd_addr_r_c[1]), .O(n12905));
    defparam rd_addr_r_0__bdd_4_lut_10965.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i6_2_lut_4_lut (.I0(\rd_addr_r[6] ), 
            .I1(rd_addr_p1_w[6]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_498[5] ), 
            .O(rd_grey_w[5]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i6_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4537_2_lut_4_lut (.I0(\rd_addr_r[6] ), .I1(rd_addr_p1_w[6]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n5920));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4537_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11520 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_6 ), 
            .I2(\REG.mem_51_6 ), .I3(rd_addr_r_c[1]), .O(n13571));
    defparam rd_addr_r_0__bdd_4_lut_11520.LUT_INIT = 16'he4aa;
    SB_LUT4 i4536_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_58_15 ), .O(n5919));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4536_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12905_bdd_4_lut (.I0(n12905), .I1(\REG.mem_9_1 ), .I2(\REG.mem_8_1 ), 
            .I3(rd_addr_r_c[1]), .O(n11302));
    defparam n12905_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4084_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_33_9 ), .O(n5467));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4084_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13571_bdd_4_lut (.I0(n13571), .I1(\REG.mem_49_6 ), .I2(\REG.mem_48_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11530));
    defparam n13571_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4535_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_58_14 ), .O(n5918));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4535_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10960 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_11 ), 
            .I2(\REG.mem_55_11 ), .I3(rd_addr_r_c[1]), .O(n12899));
    defparam rd_addr_r_0__bdd_4_lut_10960.LUT_INIT = 16'he4aa;
    SB_LUT4 i4534_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_58_13 ), .O(n5917));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4534_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4533_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_58_12 ), .O(n5916));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4533_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4532_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_58_11 ), .O(n5915));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4532_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11530 (.I0(rd_addr_r_c[2]), .I1(n13226), 
            .I2(n12836), .I3(rd_addr_r_c[3]), .O(n13565));
    defparam rd_addr_r_2__bdd_4_lut_11530.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_6__I_0_i4_3_lut (.I0(rd_addr_r_c[3]), .I1(rd_addr_p1_w[3]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_6__N_498[3] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_6__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13565_bdd_4_lut (.I0(n13565), .I1(n13418), .I2(n11500), .I3(rd_addr_r_c[3]), 
            .O(n11995));
    defparam n13565_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4531_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_58_10 ), .O(n5914));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4531_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_6__I_0_i3_3_lut (.I0(rd_addr_r_c[2]), .I1(rd_addr_p1_w[2]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_6__N_498[2] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_6__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4530_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_58_9 ), .O(n5913));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4530_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4529_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_58_8 ), .O(n5912));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4529_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4528_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_58_7 ), .O(n5911));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4528_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12899_bdd_4_lut (.I0(n12899), .I1(\REG.mem_53_11 ), .I2(\REG.mem_52_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11719));
    defparam n12899_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i88_2_lut_3_lut (.I0(n23_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n56));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i88_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i4527_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_58_6 ), .O(n5910));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4527_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4526_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_58_5 ), .O(n5909));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4526_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i87_2_lut_3_lut (.I0(n23_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n24));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i87_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i4083_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_33_8 ), .O(n5466));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4083_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10955 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_3 ), 
            .I2(\REG.mem_59_3 ), .I3(rd_addr_r_c[1]), .O(n12893));
    defparam rd_addr_r_0__bdd_4_lut_10955.LUT_INIT = 16'he4aa;
    SB_LUT4 i4525_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_58_4 ), .O(n5908));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4525_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4524_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_58_3 ), .O(n5907));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4524_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4523_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_58_2 ), .O(n5906));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4523_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12893_bdd_4_lut (.I0(n12893), .I1(\REG.mem_57_3 ), .I2(\REG.mem_56_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11125));
    defparam n12893_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_11630 (.I0(rd_addr_r_c[4]), .I1(n12554), 
            .I2(n11983), .I3(rd_addr_r_c[5]), .O(n13559));
    defparam rd_addr_r_4__bdd_4_lut_11630.LUT_INIT = 16'he4aa;
    SB_LUT4 n13559_bdd_4_lut (.I0(n13559), .I1(n13094), .I2(n11575), .I3(rd_addr_r_c[5]), 
            .O(\REG.out_raw_31__N_559 [0]));
    defparam n13559_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4522_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_58_1 ), .O(n5905));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4522_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1010_1011 (.Q(\REG.mem_10_4 ), .C(FIFO_CLK_c), .D(n5078));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4521_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_58_0 ), .O(n5904));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4521_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11515 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_3 ), 
            .I2(\REG.mem_15_3 ), .I3(rd_addr_r_c[1]), .O(n13553));
    defparam rd_addr_r_0__bdd_4_lut_11515.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i90_2_lut_3_lut_4_lut (.I0(n18_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n55));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i90_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i89_2_lut_3_lut_4_lut (.I0(n18_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n23));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i89_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_DFF i1007_1008 (.Q(\REG.mem_10_3 ), .C(FIFO_CLK_c), .D(n5077));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i120_2_lut_3_lut (.I0(n23_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n40));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i120_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i119_2_lut_3_lut (.I0(n23_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n8));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i119_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10950 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_5 ), 
            .I2(\REG.mem_35_5 ), .I3(rd_addr_r_c[1]), .O(n12887));
    defparam rd_addr_r_0__bdd_4_lut_10950.LUT_INIT = 16'he4aa;
    SB_LUT4 n13553_bdd_4_lut (.I0(n13553), .I1(\REG.mem_13_3 ), .I2(\REG.mem_12_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11056));
    defparam n13553_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12887_bdd_4_lut (.I0(n12887), .I1(\REG.mem_33_5 ), .I2(\REG.mem_32_5 ), 
            .I3(rd_addr_r_c[1]), .O(n12890));
    defparam n12887_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i23_2_lut_3_lut (.I0(n12_adj_33), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n23_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i23_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_11505 (.I0(rd_addr_r_c[4]), .I1(n11989), 
            .I2(n11995), .I3(rd_addr_r_c[5]), .O(n13547));
    defparam rd_addr_r_4__bdd_4_lut_11505.LUT_INIT = 16'he4aa;
    SB_DFF i1004_1005 (.Q(\REG.mem_10_2 ), .C(FIFO_CLK_c), .D(n5076));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1001_1002 (.Q(\REG.mem_10_1 ), .C(FIFO_CLK_c), .D(n5075));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10514 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_7 ), 
            .I2(\REG.mem_23_7 ), .I3(rd_addr_r_c[1]), .O(n12359));
    defparam rd_addr_r_0__bdd_4_lut_10514.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i40_2_lut_3_lut_4_lut (.I0(n12_adj_33), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n40_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i40_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 n13547_bdd_4_lut (.I0(n13547), .I1(n11914), .I2(n12314), .I3(rd_addr_r_c[5]), 
            .O(\REG.out_raw_31__N_559 [13]));
    defparam n13547_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i39_2_lut_3_lut_4_lut (.I0(n12_adj_33), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n39));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i39_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11060 (.I0(rd_addr_r_c[3]), .I1(n12866), 
            .I2(n11256), .I3(rd_addr_r_c[4]), .O(n12881));
    defparam rd_addr_r_3__bdd_4_lut_11060.LUT_INIT = 16'he4aa;
    SB_LUT4 n12881_bdd_4_lut (.I0(n12881), .I1(n11250), .I2(n11249), .I3(rd_addr_r_c[4]), 
            .O(n12884));
    defparam n12881_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i998_999 (.Q(\REG.mem_10_0 ), .C(FIFO_CLK_c), .D(n5074));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11500 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_6 ), 
            .I2(\REG.mem_55_6 ), .I3(rd_addr_r_c[1]), .O(n13541));
    defparam rd_addr_r_0__bdd_4_lut_11500.LUT_INIT = 16'he4aa;
    SB_LUT4 n13541_bdd_4_lut (.I0(n13541), .I1(\REG.mem_53_6 ), .I2(\REG.mem_52_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11545));
    defparam n13541_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11000 (.I0(rd_addr_r_c[1]), .I1(n11234), 
            .I2(n11235), .I3(rd_addr_r_c[2]), .O(n12875));
    defparam rd_addr_r_1__bdd_4_lut_11000.LUT_INIT = 16'he4aa;
    SB_DFF i947_948 (.Q(\REG.mem_9_15 ), .C(FIFO_CLK_c), .D(n5073));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4082_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_33_7 ), .O(n5465));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4082_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4501_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_56_15 ), .O(n5884));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4501_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4500_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_56_14 ), .O(n5883));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4500_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4499_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_56_13 ), .O(n5882));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4499_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4498_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_56_12 ), .O(n5881));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4498_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11490 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_3 ), 
            .I2(\REG.mem_19_3 ), .I3(rd_addr_r_c[1]), .O(n13535));
    defparam rd_addr_r_0__bdd_4_lut_11490.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10484 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_7 ), 
            .I2(\REG.mem_27_7 ), .I3(rd_addr_r_c[1]), .O(n12323));
    defparam rd_addr_r_0__bdd_4_lut_10484.LUT_INIT = 16'he4aa;
    SB_DFF i944_945 (.Q(\REG.mem_9_14 ), .C(FIFO_CLK_c), .D(n5072));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12875_bdd_4_lut (.I0(n12875), .I1(n11226), .I2(n11225), .I3(rd_addr_r_c[2]), 
            .O(n12878));
    defparam n12875_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4497_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_56_11 ), .O(n5880));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4497_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13535_bdd_4_lut (.I0(n13535), .I1(\REG.mem_17_3 ), .I2(\REG.mem_16_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11059));
    defparam n13535_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i20_2_lut (.I0(n11), .I1(wr_addr_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n20_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i20_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4496_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_56_10 ), .O(n5879));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4496_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i146_147 (.Q(\REG.mem_1_4 ), .C(FIFO_CLK_c), .D(n4837));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4495_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_56_9 ), .O(n5878));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4495_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10935 (.I0(rd_addr_r_c[1]), .I1(n11213), 
            .I2(n11214), .I3(rd_addr_r_c[2]), .O(n12869));
    defparam rd_addr_r_1__bdd_4_lut_10935.LUT_INIT = 16'he4aa;
    SB_LUT4 i4494_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_56_8 ), .O(n5877));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4494_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4493_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_56_7 ), .O(n5876));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4493_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4492_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_56_6 ), .O(n5875));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4492_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i941_942 (.Q(\REG.mem_9_13 ), .C(FIFO_CLK_c), .D(n5071));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11525 (.I0(rd_addr_r_c[3]), .I1(n12722), 
            .I2(n11052), .I3(rd_addr_r_c[4]), .O(n13529));
    defparam rd_addr_r_3__bdd_4_lut_11525.LUT_INIT = 16'he4aa;
    SB_DFF i938_939 (.Q(\REG.mem_9_12 ), .C(FIFO_CLK_c), .D(n5070));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4491_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_56_5 ), .O(n5874));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4491_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9672_3_lut (.I0(\REG.mem_56_7 ), .I1(\REG.mem_57_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11510));
    defparam i9672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12359_bdd_4_lut (.I0(n12359), .I1(\REG.mem_21_7 ), .I2(\REG.mem_20_7 ), 
            .I3(rd_addr_r_c[1]), .O(n12362));
    defparam n12359_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12869_bdd_4_lut (.I0(n12869), .I1(n11208), .I2(n11207), .I3(rd_addr_r_c[2]), 
            .O(n12872));
    defparam n12869_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9673_3_lut (.I0(\REG.mem_58_7 ), .I1(\REG.mem_59_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11511));
    defparam i9673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10930 (.I0(rd_addr_r_c[1]), .I1(n11189), 
            .I2(n11190), .I3(rd_addr_r_c[2]), .O(n12863));
    defparam rd_addr_r_1__bdd_4_lut_10930.LUT_INIT = 16'he4aa;
    SB_DFF i935_936 (.Q(\REG.mem_9_11 ), .C(FIFO_CLK_c), .D(n5069));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4490_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_56_4 ), .O(n5873));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4490_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12863_bdd_4_lut (.I0(n12863), .I1(n11178), .I2(n11177), .I3(rd_addr_r_c[2]), 
            .O(n12866));
    defparam n12863_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4489_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_56_3 ), .O(n5872));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4489_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4488_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_56_2 ), .O(n5871));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4488_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4487_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_56_1 ), .O(n5870));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4487_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_33 (.I0(DEBUG_3_c), .I1(get_next_word), .I2(GND_net), 
            .I3(GND_net), .O(rd_fifo_en_w));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i1_2_lut_adj_33.LUT_INIT = 16'h4444;
    SB_LUT4 n13529_bdd_4_lut (.I0(n13529), .I1(n11028), .I2(n11027), .I3(rd_addr_r_c[4]), 
            .O(n13532));
    defparam n13529_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4482_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_56_0 ), .O(n5865));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4482_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10509 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_15 ), 
            .I2(\REG.mem_47_15 ), .I3(rd_addr_r_c[1]), .O(n12353));
    defparam rd_addr_r_0__bdd_4_lut_10509.LUT_INIT = 16'he4aa;
    SB_DFF i149_150 (.Q(\REG.mem_1_5 ), .C(FIFO_CLK_c), .D(n4835));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i932_933 (.Q(\REG.mem_9_10 ), .C(FIFO_CLK_c), .D(n5068));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i929_930 (.Q(\REG.mem_9_9 ), .C(FIFO_CLK_c), .D(n5067));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10945 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_11 ), 
            .I2(\REG.mem_59_11 ), .I3(rd_addr_r_c[1]), .O(n12857));
    defparam rd_addr_r_0__bdd_4_lut_10945.LUT_INIT = 16'he4aa;
    SB_LUT4 n12857_bdd_4_lut (.I0(n12857), .I1(\REG.mem_57_11 ), .I2(\REG.mem_56_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11722));
    defparam n12857_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i926_927 (.Q(\REG.mem_9_8 ), .C(FIFO_CLK_c), .D(n5066));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9694_3_lut (.I0(\REG.mem_62_7 ), .I1(\REG.mem_63_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11532));
    defparam i9694_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i923_924 (.Q(\REG.mem_9_7 ), .C(FIFO_CLK_c), .D(n5065));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11535 (.I0(rd_addr_r_c[1]), .I1(n11435), 
            .I2(n11436), .I3(rd_addr_r_c[2]), .O(n13523));
    defparam rd_addr_r_1__bdd_4_lut_11535.LUT_INIT = 16'he4aa;
    SB_LUT4 n13523_bdd_4_lut (.I0(n13523), .I1(n11427), .I2(n11426), .I3(rd_addr_r_c[2]), 
            .O(n11550));
    defparam n13523_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9693_3_lut (.I0(\REG.mem_60_7 ), .I1(\REG.mem_61_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11531));
    defparam i9693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i53_2_lut_3_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n53_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i53_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i86_2_lut_3_lut_4_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n57));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i86_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11485 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_3 ), 
            .I2(\REG.mem_23_3 ), .I3(rd_addr_r_c[1]), .O(n13517));
    defparam rd_addr_r_0__bdd_4_lut_11485.LUT_INIT = 16'he4aa;
    SB_DFF i920_921 (.Q(\REG.mem_9_6 ), .C(FIFO_CLK_c), .D(n5064));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13517_bdd_4_lut (.I0(n13517), .I1(\REG.mem_21_3 ), .I2(\REG.mem_20_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11065));
    defparam n13517_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i85_2_lut_3_lut_4_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n25));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i85_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i4081_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_33_6 ), .O(n5464));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4081_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11470 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_14 ), 
            .I2(\REG.mem_51_14 ), .I3(rd_addr_r_c[1]), .O(n13511));
    defparam rd_addr_r_0__bdd_4_lut_11470.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i2_2_lut_4_lut (.I0(rd_addr_r_c[1]), 
            .I1(rd_addr_p1_w[1]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_498[2] ), 
            .O(rd_grey_w[1]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i2_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 n13511_bdd_4_lut (.I0(n13511), .I1(\REG.mem_49_14 ), .I2(\REG.mem_48_14 ), 
            .I3(rd_addr_r_c[1]), .O(n12010));
    defparam n13511_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i917_918 (.Q(\REG.mem_9_5 ), .C(FIFO_CLK_c), .D(n5063));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10920 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_0 ), 
            .I2(\REG.mem_23_0 ), .I3(rd_addr_r_c[1]), .O(n12851));
    defparam rd_addr_r_0__bdd_4_lut_10920.LUT_INIT = 16'he4aa;
    SB_LUT4 n12851_bdd_4_lut (.I0(n12851), .I1(\REG.mem_21_0 ), .I2(\REG.mem_20_0 ), 
            .I3(rd_addr_r_c[1]), .O(n12854));
    defparam n12851_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11465 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_14 ), 
            .I2(\REG.mem_55_14 ), .I3(rd_addr_r_c[1]), .O(n13505));
    defparam rd_addr_r_0__bdd_4_lut_11465.LUT_INIT = 16'he4aa;
    SB_LUT4 i4542_2_lut_4_lut (.I0(rd_addr_r_c[1]), .I1(rd_addr_p1_w[1]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n5925));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4542_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 n13505_bdd_4_lut (.I0(n13505), .I1(\REG.mem_53_14 ), .I2(\REG.mem_52_14 ), 
            .I3(rd_addr_r_c[1]), .O(n12016));
    defparam n13505_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i914_915 (.Q(\REG.mem_9_4 ), .C(FIFO_CLK_c), .D(n5062));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4080_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_33_5 ), .O(n5463));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4080_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_34 (.I0(rp_sync2_r[5]), .I1(rp_sync2_r[4]), .I2(rp_sync2_r[6]), 
            .I3(GND_net), .O(rp_sync_w[4]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i2_3_lut_adj_34.LUT_INIT = 16'h6969;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i1_2_lut_4_lut (.I0(rd_addr_r_c[1]), 
            .I1(rd_addr_p1_w[1]), .I2(rd_fifo_en_w), .I3(rd_addr_nxt_c_6__N_498[0]), 
            .O(rd_grey_w[0]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i1_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i1_2_lut_adj_35 (.I0(rp_sync2_r[3]), .I1(rp_sync_w[4]), .I2(GND_net), 
            .I3(GND_net), .O(rp_sync_w[3]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_adj_35.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_36 (.I0(rp_sync2_r[1]), .I1(rp_sync_w[2]), .I2(GND_net), 
            .I3(GND_net), .O(rp_sync_w[1]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_adj_36.LUT_INIT = 16'h6666;
    SB_LUT4 i3483_2_lut_4_lut (.I0(wr_addr_r[0]), .I1(wr_addr_p1_w[0]), 
            .I2(wr_sig_mv_w), .I3(reset_per_frame), .O(n4866));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i3483_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 rp_sync2_r_6__I_0_136_i1_2_lut (.I0(rp_sync2_r[5]), .I1(rp_sync2_r[6]), 
            .I2(GND_net), .I3(GND_net), .O(rp_sync_w[5]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam rp_sync2_r_6__I_0_136_i1_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i1_2_lut_4_lut (.I0(wr_addr_r[0]), .I1(wr_addr_p1_w[0]), 
            .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[1] ), .O(wr_grey_w[0]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i1_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_DFF i911_912 (.Q(\REG.mem_9_3 ), .C(FIFO_CLK_c), .D(n5061));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3561_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_0_0 ), .O(n4944));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3561_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3541_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_0_15 ), .O(n4924));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3541_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3542_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_0_14 ), .O(n4925));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3542_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3543_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_0_13 ), .O(n4926));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3543_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3544_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_0_12 ), .O(n4927));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3544_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3545_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_0_11 ), .O(n4928));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3545_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i908_909 (.Q(\REG.mem_9_2 ), .C(FIFO_CLK_c), .D(n5060));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i905_906 (.Q(\REG.mem_9_1 ), .C(FIFO_CLK_c), .D(n5059));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i902_903 (.Q(\REG.mem_9_0 ), .C(FIFO_CLK_c), .D(n5057));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i851_852 (.Q(\REG.mem_8_15 ), .C(FIFO_CLK_c), .D(n5056));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i848_849 (.Q(\REG.mem_8_14 ), .C(FIFO_CLK_c), .D(n5055));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i845_846 (.Q(\REG.mem_8_13 ), .C(FIFO_CLK_c), .D(n5054));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i842_843 (.Q(\REG.mem_8_12 ), .C(FIFO_CLK_c), .D(n5053));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i839_840 (.Q(\REG.mem_8_11 ), .C(FIFO_CLK_c), .D(n5052));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i836_837 (.Q(\REG.mem_8_10 ), .C(FIFO_CLK_c), .D(n5051));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i833_834 (.Q(\REG.mem_8_9 ), .C(FIFO_CLK_c), .D(n5050));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i830_831 (.Q(\REG.mem_8_8 ), .C(FIFO_CLK_c), .D(n5049));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i827_828 (.Q(\REG.mem_8_7 ), .C(FIFO_CLK_c), .D(n5048));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i824_825 (.Q(\REG.mem_8_6 ), .C(FIFO_CLK_c), .D(n5047));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i821_822 (.Q(\REG.mem_8_5 ), .C(FIFO_CLK_c), .D(n5046));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i818_819 (.Q(\REG.mem_8_4 ), .C(FIFO_CLK_c), .D(n5045));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i815_816 (.Q(\REG.mem_8_3 ), .C(FIFO_CLK_c), .D(n5044));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i812_813 (.Q(\REG.mem_8_2 ), .C(FIFO_CLK_c), .D(n5043));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i809_810 (.Q(\REG.mem_8_1 ), .C(FIFO_CLK_c), .D(n5042));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i806_807 (.Q(\REG.mem_8_0 ), .C(FIFO_CLK_c), .D(n5041));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i755_756 (.Q(\REG.mem_7_15 ), .C(FIFO_CLK_c), .D(n5040));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i752_753 (.Q(\REG.mem_7_14 ), .C(FIFO_CLK_c), .D(n5039));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i749_750 (.Q(\REG.mem_7_13 ), .C(FIFO_CLK_c), .D(n5038));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i746_747 (.Q(\REG.mem_7_12 ), .C(FIFO_CLK_c), .D(n5037));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i743_744 (.Q(\REG.mem_7_11 ), .C(FIFO_CLK_c), .D(n5036));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i740_741 (.Q(\REG.mem_7_10 ), .C(FIFO_CLK_c), .D(n5035));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i737_738 (.Q(\REG.mem_7_9 ), .C(FIFO_CLK_c), .D(n5034));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i734_735 (.Q(\REG.mem_7_8 ), .C(FIFO_CLK_c), .D(n5033));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i731_732 (.Q(\REG.mem_7_7 ), .C(FIFO_CLK_c), .D(n5032));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i728_729 (.Q(\REG.mem_7_6 ), .C(FIFO_CLK_c), .D(n5031));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i725_726 (.Q(\REG.mem_7_5 ), .C(FIFO_CLK_c), .D(n5030));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i722_723 (.Q(\REG.mem_7_4 ), .C(FIFO_CLK_c), .D(n5029));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i719_720 (.Q(\REG.mem_7_3 ), .C(FIFO_CLK_c), .D(n5028));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i716_717 (.Q(\REG.mem_7_2 ), .C(FIFO_CLK_c), .D(n5027));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i713_714 (.Q(\REG.mem_7_1 ), .C(FIFO_CLK_c), .D(n5026));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i710_711 (.Q(\REG.mem_7_0 ), .C(FIFO_CLK_c), .D(n5025));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i659_660 (.Q(\REG.mem_6_15 ), .C(FIFO_CLK_c), .D(n5024));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i656_657 (.Q(\REG.mem_6_14 ), .C(FIFO_CLK_c), .D(n5023));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i653_654 (.Q(\REG.mem_6_13 ), .C(FIFO_CLK_c), .D(n5022));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i650_651 (.Q(\REG.mem_6_12 ), .C(FIFO_CLK_c), .D(n5021));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i647_648 (.Q(\REG.mem_6_11 ), .C(FIFO_CLK_c), .D(n5020));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i644_645 (.Q(\REG.mem_6_10 ), .C(FIFO_CLK_c), .D(n5019));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i641_642 (.Q(\REG.mem_6_9 ), .C(FIFO_CLK_c), .D(n5018));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i638_639 (.Q(\REG.mem_6_8 ), .C(FIFO_CLK_c), .D(n5017));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i635_636 (.Q(\REG.mem_6_7 ), .C(FIFO_CLK_c), .D(n5016));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i632_633 (.Q(\REG.mem_6_6 ), .C(FIFO_CLK_c), .D(n5015));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i629_630 (.Q(\REG.mem_6_5 ), .C(FIFO_CLK_c), .D(n5014));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i626_627 (.Q(\REG.mem_6_4 ), .C(FIFO_CLK_c), .D(n5013));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i623_624 (.Q(\REG.mem_6_3 ), .C(FIFO_CLK_c), .D(n5012));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i620_621 (.Q(\REG.mem_6_2 ), .C(FIFO_CLK_c), .D(n5011));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i617_618 (.Q(\REG.mem_6_1 ), .C(FIFO_CLK_c), .D(n5010));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i614_615 (.Q(\REG.mem_6_0 ), .C(FIFO_CLK_c), .D(n5009));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i563_564 (.Q(\REG.mem_5_15 ), .C(FIFO_CLK_c), .D(n5008));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i560_561 (.Q(\REG.mem_5_14 ), .C(FIFO_CLK_c), .D(n5007));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i557_558 (.Q(\REG.mem_5_13 ), .C(FIFO_CLK_c), .D(n5006));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i554_555 (.Q(\REG.mem_5_12 ), .C(FIFO_CLK_c), .D(n5005));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i551_552 (.Q(\REG.mem_5_11 ), .C(FIFO_CLK_c), .D(n5004));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i548_549 (.Q(\REG.mem_5_10 ), .C(FIFO_CLK_c), .D(n5003));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i545_546 (.Q(\REG.mem_5_9 ), .C(FIFO_CLK_c), .D(n5002));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i542_543 (.Q(\REG.mem_5_8 ), .C(FIFO_CLK_c), .D(n5001));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i539_540 (.Q(\REG.mem_5_7 ), .C(FIFO_CLK_c), .D(n5000));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i536_537 (.Q(\REG.mem_5_6 ), .C(FIFO_CLK_c), .D(n4999));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i533_534 (.Q(\REG.mem_5_5 ), .C(FIFO_CLK_c), .D(n4998));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i530_531 (.Q(\REG.mem_5_4 ), .C(FIFO_CLK_c), .D(n4997));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i527_528 (.Q(\REG.mem_5_3 ), .C(FIFO_CLK_c), .D(n4996));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i524_525 (.Q(\REG.mem_5_2 ), .C(FIFO_CLK_c), .D(n4995));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i521_522 (.Q(\REG.mem_5_1 ), .C(FIFO_CLK_c), .D(n4994));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i518_519 (.Q(\REG.mem_5_0 ), .C(FIFO_CLK_c), .D(n4993));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i467_468 (.Q(\REG.mem_4_15 ), .C(FIFO_CLK_c), .D(n4992));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i464_465 (.Q(\REG.mem_4_14 ), .C(FIFO_CLK_c), .D(n4991));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i461_462 (.Q(\REG.mem_4_13 ), .C(FIFO_CLK_c), .D(n4990));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i458_459 (.Q(\REG.mem_4_12 ), .C(FIFO_CLK_c), .D(n4989));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i455_456 (.Q(\REG.mem_4_11 ), .C(FIFO_CLK_c), .D(n4988));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i452_453 (.Q(\REG.mem_4_10 ), .C(FIFO_CLK_c), .D(n4987));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i449_450 (.Q(\REG.mem_4_9 ), .C(FIFO_CLK_c), .D(n4986));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i446_447 (.Q(\REG.mem_4_8 ), .C(FIFO_CLK_c), .D(n4985));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i443_444 (.Q(\REG.mem_4_7 ), .C(FIFO_CLK_c), .D(n4984));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i440_441 (.Q(\REG.mem_4_6 ), .C(FIFO_CLK_c), .D(n4983));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i437_438 (.Q(\REG.mem_4_5 ), .C(FIFO_CLK_c), .D(n4982));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i434_435 (.Q(\REG.mem_4_4 ), .C(FIFO_CLK_c), .D(n4981));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i431_432 (.Q(\REG.mem_4_3 ), .C(FIFO_CLK_c), .D(n4980));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i428_429 (.Q(\REG.mem_4_2 ), .C(FIFO_CLK_c), .D(n4979));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i425_426 (.Q(\REG.mem_4_1 ), .C(FIFO_CLK_c), .D(n4978));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i422_423 (.Q(\REG.mem_4_0 ), .C(FIFO_CLK_c), .D(n4977));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i371_372 (.Q(\REG.mem_3_15 ), .C(FIFO_CLK_c), .D(n4976));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i368_369 (.Q(\REG.mem_3_14 ), .C(FIFO_CLK_c), .D(n4975));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i365_366 (.Q(\REG.mem_3_13 ), .C(FIFO_CLK_c), .D(n4974));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i362_363 (.Q(\REG.mem_3_12 ), .C(FIFO_CLK_c), .D(n4973));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i359_360 (.Q(\REG.mem_3_11 ), .C(FIFO_CLK_c), .D(n4972));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i356_357 (.Q(\REG.mem_3_10 ), .C(FIFO_CLK_c), .D(n4971));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i353_354 (.Q(\REG.mem_3_9 ), .C(FIFO_CLK_c), .D(n4970));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i350_351 (.Q(\REG.mem_3_8 ), .C(FIFO_CLK_c), .D(n4969));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12317_bdd_4_lut (.I0(n12317), .I1(n11143), .I2(n11122), .I3(rd_addr_r_c[3]), 
            .O(n12320));
    defparam n12317_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12353_bdd_4_lut (.I0(n12353), .I1(\REG.mem_45_15 ), .I2(\REG.mem_44_15 ), 
            .I3(rd_addr_r_c[1]), .O(n12356));
    defparam n12353_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3546_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_0_10 ), .O(n4929));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3546_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3547_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_0_9 ), .O(n4930));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3547_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11475 (.I0(rd_addr_r_c[1]), .I1(n11468), 
            .I2(n11469), .I3(rd_addr_r_c[2]), .O(n13499));
    defparam rd_addr_r_1__bdd_4_lut_11475.LUT_INIT = 16'he4aa;
    SB_LUT4 i9009_4_lut (.I0(wr_addr_r[1]), .I1(wr_addr_r[3]), .I2(rp_sync_w[1]), 
            .I3(rp_sync_w[3]), .O(n10845));
    defparam i9009_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 n13499_bdd_4_lut (.I0(n13499), .I1(n11457), .I2(n11456), .I3(rd_addr_r_c[2]), 
            .O(n11559));
    defparam n13499_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_p1_w_6__I_0_2_lut (.I0(wr_addr_p1_w[6]), .I1(rp_sync2_r[6]), 
            .I2(GND_net), .I3(GND_net), .O(full_max_w));   // src/fifo_dc_32_lut_gen.v(296[27:88])
    defparam wr_addr_p1_w_6__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10915 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_3 ), 
            .I2(\REG.mem_63_3 ), .I3(rd_addr_r_c[1]), .O(n12845));
    defparam rd_addr_r_0__bdd_4_lut_10915.LUT_INIT = 16'he4aa;
    SB_LUT4 i9013_4_lut (.I0(wr_addr_p1_w[4]), .I1(wr_addr_p1_w[1]), .I2(rp_sync_w[4]), 
            .I3(rp_sync_w[1]), .O(n10849));
    defparam i9013_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 i9045_4_lut (.I0(wr_addr_p1_w[5]), .I1(wr_addr_p1_w[3]), .I2(rp_sync_w[5]), 
            .I3(rp_sync_w[3]), .O(n10881));
    defparam i9045_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 i5_4_lut_adj_37 (.I0(wr_addr_p1_w[0]), .I1(n10849), .I2(full_max_w), 
            .I3(rp_sync_w[0]), .O(n12_adj_35));
    defparam i5_4_lut_adj_37.LUT_INIT = 16'h1020;
    SB_LUT4 wr_addr_r_5__I_0_i3_2_lut (.I0(wr_addr_r[2]), .I1(rp_sync_w[2]), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_36));   // src/fifo_dc_32_lut_gen.v(295[31:67])
    defparam wr_addr_r_5__I_0_i3_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i9110_4_lut (.I0(wr_addr_r[0]), .I1(n10845), .I2(n6_adj_37), 
            .I3(rp_sync_w[0]), .O(n10947));
    defparam i9110_4_lut.LUT_INIT = 16'hfefd;
    SB_LUT4 i10355_4_lut (.I0(wr_addr_p1_w[2]), .I1(n12_adj_35), .I2(n10881), 
            .I3(rp_sync_w[2]), .O(n12032));   // src/fifo_dc_32_lut_gen.v(300[45:114])
    defparam i10355_4_lut.LUT_INIT = 16'h0408;
    SB_LUT4 i10354_4_lut (.I0(wr_addr_r[4]), .I1(full_o), .I2(rp_sync_w[4]), 
            .I3(n3_adj_36), .O(n12033));   // src/fifo_dc_32_lut_gen.v(300[45:114])
    defparam i10354_4_lut.LUT_INIT = 16'h0048;
    SB_LUT4 full_nxt_c_I_6_4_lut (.I0(n12033), .I1(n12032), .I2(wr_sig_mv_w), 
            .I3(n10947), .O(full_nxt_c_N_626));   // src/fifo_dc_32_lut_gen.v(300[45:114])
    defparam full_nxt_c_I_6_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i1_2_lut_adj_38 (.I0(dc32_fifo_almost_full), .I1(DEBUG_1_c_c), 
            .I2(GND_net), .I3(GND_net), .O(FT_OE_N_420));   // src/fifo_dc_32_lut_gen.v(410[29] 422[32])
    defparam i1_2_lut_adj_38.LUT_INIT = 16'heeee;
    SB_LUT4 n12845_bdd_4_lut (.I0(n12845), .I1(\REG.mem_61_3 ), .I2(\REG.mem_60_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11128));
    defparam n12845_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3548_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_0_8 ), .O(n4931));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3548_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11455 (.I0(rd_addr_r_c[1]), .I1(n11507), 
            .I2(n11508), .I3(rd_addr_r_c[2]), .O(n13493));
    defparam rd_addr_r_1__bdd_4_lut_11455.LUT_INIT = 16'he4aa;
    SB_LUT4 n13493_bdd_4_lut (.I0(n13493), .I1(n11496), .I2(n11495), .I3(rd_addr_r_c[2]), 
            .O(n11562));
    defparam n13493_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i161_162 (.Q(\REG.mem_1_9 ), .C(FIFO_CLK_c), .D(n4833));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11460 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_8 ), 
            .I2(\REG.mem_3_8 ), .I3(rd_addr_r_c[1]), .O(n13487));
    defparam rd_addr_r_0__bdd_4_lut_11460.LUT_INIT = 16'he4aa;
    SB_LUT4 n13487_bdd_4_lut (.I0(n13487), .I1(\REG.mem_1_8 ), .I2(\REG.mem_0_8 ), 
            .I3(rd_addr_r_c[1]), .O(n13490));
    defparam n13487_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10940 (.I0(rd_addr_r_c[3]), .I1(n12746), 
            .I2(n11070), .I3(rd_addr_r_c[4]), .O(n12839));
    defparam rd_addr_r_3__bdd_4_lut_10940.LUT_INIT = 16'he4aa;
    SB_LUT4 i3549_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_0_7 ), .O(n4932));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3549_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11480 (.I0(rd_addr_r_c[3]), .I1(n11888), 
            .I2(n11889), .I3(rd_addr_r_c[4]), .O(n13481));
    defparam rd_addr_r_3__bdd_4_lut_11480.LUT_INIT = 16'he4aa;
    SB_LUT4 n13481_bdd_4_lut (.I0(n13481), .I1(n11877), .I2(n13394), .I3(rd_addr_r_c[4]), 
            .O(n13484));
    defparam n13481_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i179_180 (.Q(\REG.mem_1_15 ), .C(FIFO_CLK_c), .D(n4832));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12839_bdd_4_lut (.I0(n12839), .I1(n11025), .I2(n12692), .I3(rd_addr_r_c[4]), 
            .O(n12842));
    defparam n12839_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_en_i_I_0_2_lut (.I0(DEBUG_5_c), .I1(full_o), .I2(GND_net), 
            .I3(GND_net), .O(wr_sig_mv_w));   // src/fifo_dc_32_lut_gen.v(293[28:49])
    defparam wr_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10910 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_13 ), 
            .I2(\REG.mem_63_13 ), .I3(rd_addr_r_c[1]), .O(n12833));
    defparam rd_addr_r_0__bdd_4_lut_10910.LUT_INIT = 16'he4aa;
    SB_LUT4 n12833_bdd_4_lut (.I0(n12833), .I1(\REG.mem_61_13 ), .I2(\REG.mem_60_13 ), 
            .I3(rd_addr_r_c[1]), .O(n12836));
    defparam n12833_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11445 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_3 ), 
            .I2(\REG.mem_27_3 ), .I3(rd_addr_r_c[1]), .O(n13475));
    defparam rd_addr_r_0__bdd_4_lut_11445.LUT_INIT = 16'he4aa;
    SB_DFF i164_165 (.Q(\REG.mem_1_10 ), .C(FIFO_CLK_c), .D(n4831));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3550_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_0_6 ), .O(n4933));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3550_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i18_2_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n18_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i18_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3551_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_0_5 ), .O(n4934));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3551_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3552_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_0_4 ), .O(n4935));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3552_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13475_bdd_4_lut (.I0(n13475), .I1(\REG.mem_25_3 ), .I2(\REG.mem_24_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11068));
    defparam n13475_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3557_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_0_3 ), .O(n4940));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3557_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10900 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_0 ), 
            .I2(\REG.mem_27_0 ), .I3(rd_addr_r_c[1]), .O(n12827));
    defparam rd_addr_r_0__bdd_4_lut_10900.LUT_INIT = 16'he4aa;
    SB_LUT4 i3558_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_0_2 ), .O(n4941));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3558_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12827_bdd_4_lut (.I0(n12827), .I1(\REG.mem_25_0 ), .I2(\REG.mem_24_0 ), 
            .I3(rd_addr_r_c[1]), .O(n12830));
    defparam n12827_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3560_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_0_1 ), .O(n4943));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3560_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11435 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_5 ), 
            .I2(\REG.mem_11_5 ), .I3(rd_addr_r_c[1]), .O(n13469));
    defparam rd_addr_r_0__bdd_4_lut_11435.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i38_2_lut_3_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n38));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i38_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10895 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_9 ), 
            .I2(\REG.mem_47_9 ), .I3(rd_addr_r_c[1]), .O(n12821));
    defparam rd_addr_r_0__bdd_4_lut_10895.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i102_2_lut_3_lut_4_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n49));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i102_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 n13469_bdd_4_lut (.I0(n13469), .I1(\REG.mem_9_5 ), .I2(\REG.mem_8_5 ), 
            .I3(rd_addr_r_c[1]), .O(n13472));
    defparam n13469_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12821_bdd_4_lut (.I0(n12821), .I1(\REG.mem_45_9 ), .I2(\REG.mem_44_9 ), 
            .I3(rd_addr_r_c[1]), .O(n12824));
    defparam n12821_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i101_2_lut_3_lut_4_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n17));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i101_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i116_2_lut_3_lut (.I0(n36), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n42));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i116_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i115_2_lut_3_lut (.I0(n36), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n10));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i115_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10990 (.I0(rd_addr_r_c[2]), .I1(n11464), 
            .I2(n11485), .I3(rd_addr_r_c[3]), .O(n12815));
    defparam rd_addr_r_2__bdd_4_lut_10990.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11450 (.I0(rd_addr_r_c[1]), .I1(n11915), 
            .I2(n11916), .I3(rd_addr_r_c[2]), .O(n13463));
    defparam rd_addr_r_1__bdd_4_lut_11450.LUT_INIT = 16'he4aa;
    SB_LUT4 i4079_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_33_4 ), .O(n5462));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4079_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13463_bdd_4_lut (.I0(n13463), .I1(n11892), .I2(n11891), .I3(rd_addr_r_c[2]), 
            .O(n11070));
    defparam n13463_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10504 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_2 ), 
            .I2(\REG.mem_15_2 ), .I3(rd_addr_r_c[1]), .O(n12347));
    defparam rd_addr_r_0__bdd_4_lut_10504.LUT_INIT = 16'he4aa;
    SB_LUT4 n12815_bdd_4_lut (.I0(n12815), .I1(n11407), .I2(n12374), .I3(rd_addr_r_c[3]), 
            .O(n11728));
    defparam n12815_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10890 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_1 ), 
            .I2(\REG.mem_63_1 ), .I3(rd_addr_r_c[1]), .O(n12809));
    defparam rd_addr_r_0__bdd_4_lut_10890.LUT_INIT = 16'he4aa;
    SB_LUT4 n12809_bdd_4_lut (.I0(n12809), .I1(\REG.mem_61_1 ), .I2(\REG.mem_60_1 ), 
            .I3(rd_addr_r_c[1]), .O(n12812));
    defparam n12809_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4078_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_33_3 ), .O(n5461));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4078_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11430 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_12 ), 
            .I2(\REG.mem_11_12 ), .I3(rd_addr_r_c[1]), .O(n13457));
    defparam rd_addr_r_0__bdd_4_lut_11430.LUT_INIT = 16'he4aa;
    SB_LUT4 n13457_bdd_4_lut (.I0(n13457), .I1(\REG.mem_9_12 ), .I2(\REG.mem_8_12 ), 
            .I3(rd_addr_r_c[1]), .O(n13460));
    defparam n13457_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i347_348 (.Q(\REG.mem_3_7 ), .C(FIFO_CLK_c), .D(n4968));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i344_345 (.Q(\REG.mem_3_6 ), .C(FIFO_CLK_c), .D(n4967));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9409_3_lut (.I0(\REG.mem_30_9 ), .I1(\REG.mem_31_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11247));
    defparam i9409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9408_3_lut (.I0(\REG.mem_28_9 ), .I1(\REG.mem_29_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11246));
    defparam i9408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i15_2_lut (.I0(n12_adj_33), .I1(wr_addr_r[2]), 
            .I2(GND_net), .I3(GND_net), .O(n15_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i15_2_lut.LUT_INIT = 16'h8888;
    SB_DFF i341_342 (.Q(\REG.mem_3_5 ), .C(FIFO_CLK_c), .D(n4966));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i338_339 (.Q(\REG.mem_3_4 ), .C(FIFO_CLK_c), .D(n4965));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i132_2_lut_3_lut (.I0(n35), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n34));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i132_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i335_336 (.Q(\REG.mem_3_3 ), .C(FIFO_CLK_c), .D(n4964));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11425 (.I0(rd_addr_r_c[1]), .I1(n12026), 
            .I2(n12027), .I3(rd_addr_r_c[2]), .O(n13451));
    defparam rd_addr_r_1__bdd_4_lut_11425.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10925 (.I0(rd_addr_r_c[1]), .I1(n11984), 
            .I2(n11985), .I3(rd_addr_r_c[2]), .O(n12797));
    defparam rd_addr_r_1__bdd_4_lut_10925.LUT_INIT = 16'he4aa;
    SB_LUT4 i4452_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_54_15 ), .O(n5835));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4452_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13451_bdd_4_lut (.I0(n13451), .I1(n11973), .I2(n11972), .I3(rd_addr_r_c[2]), 
            .O(n13454));
    defparam n13451_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4451_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_54_14 ), .O(n5834));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4451_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12797_bdd_4_lut (.I0(n12797), .I1(n11979), .I2(n11978), .I3(rd_addr_r_c[2]), 
            .O(n12800));
    defparam n12797_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4450_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_54_13 ), .O(n5833));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4450_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4449_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_54_12 ), .O(n5832));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4449_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4448_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_54_11 ), .O(n5831));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4448_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11420 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_8 ), 
            .I2(\REG.mem_31_8 ), .I3(rd_addr_r_c[1]), .O(n13445));
    defparam rd_addr_r_0__bdd_4_lut_11420.LUT_INIT = 16'he4aa;
    SB_LUT4 n13445_bdd_4_lut (.I0(n13445), .I1(\REG.mem_29_8 ), .I2(\REG.mem_28_8 ), 
            .I3(rd_addr_r_c[1]), .O(n13448));
    defparam n13445_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i332_333 (.Q(\REG.mem_3_2 ), .C(FIFO_CLK_c), .D(n4963));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4447_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_54_10 ), .O(n5830));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4447_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4446_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_54_9 ), .O(n5829));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4446_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4445_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_54_8 ), .O(n5828));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4445_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4077_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_33_2 ), .O(n5460));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4077_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i131_2_lut_3_lut (.I0(n35), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n2));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i131_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i4444_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_54_7 ), .O(n5827));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4444_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4443_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_54_6 ), .O(n5826));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4443_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4442_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_54_5 ), .O(n5825));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4442_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10885 (.I0(rd_addr_r_c[2]), .I1(n11044), 
            .I2(n11056), .I3(rd_addr_r_c[3]), .O(n12791));
    defparam rd_addr_r_2__bdd_4_lut_10885.LUT_INIT = 16'he4aa;
    SB_LUT4 n12791_bdd_4_lut (.I0(n12791), .I1(n11041), .I2(n11035), .I3(rd_addr_r_c[3]), 
            .O(n11131));
    defparam n12791_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4441_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_54_4 ), .O(n5824));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4441_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11410 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_1 ), 
            .I2(\REG.mem_43_1 ), .I3(rd_addr_r_c[1]), .O(n13439));
    defparam rd_addr_r_0__bdd_4_lut_11410.LUT_INIT = 16'he4aa;
    SB_LUT4 i4440_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_54_3 ), .O(n5823));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4440_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10905 (.I0(rd_addr_r_c[3]), .I1(n12020), 
            .I2(n12021), .I3(rd_addr_r_c[4]), .O(n12785));
    defparam rd_addr_r_3__bdd_4_lut_10905.LUT_INIT = 16'he4aa;
    SB_LUT4 n13439_bdd_4_lut (.I0(n13439), .I1(\REG.mem_41_1 ), .I2(\REG.mem_40_1 ), 
            .I3(rd_addr_r_c[1]), .O(n13442));
    defparam n13439_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i329_330 (.Q(\REG.mem_3_1 ), .C(FIFO_CLK_c), .D(n4962));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4439_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_54_2 ), .O(n5822));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4439_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12785_bdd_4_lut (.I0(n12785), .I1(n12003), .I2(n12002), .I3(rd_addr_r_c[4]), 
            .O(n12788));
    defparam n12785_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i326_327 (.Q(\REG.mem_3_0 ), .C(FIFO_CLK_c), .D(n4961));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12347_bdd_4_lut (.I0(n12347), .I1(\REG.mem_13_2 ), .I2(\REG.mem_12_2 ), 
            .I3(rd_addr_r_c[1]), .O(n12350));
    defparam n12347_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10880 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_12 ), 
            .I2(\REG.mem_47_12 ), .I3(rd_addr_r_c[1]), .O(n12779));
    defparam rd_addr_r_0__bdd_4_lut_10880.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i36_2_lut_3_lut (.I0(n11), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n36));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i36_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i4438_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_54_1 ), .O(n5821));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4438_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4437_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_54_0 ), .O(n5820));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4437_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i275_276 (.Q(\REG.mem_2_15 ), .C(FIFO_CLK_c), .D(n4960));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11415 (.I0(rd_addr_r_c[1]), .I1(n11465), 
            .I2(n11466), .I3(rd_addr_r_c[2]), .O(n13433));
    defparam rd_addr_r_1__bdd_4_lut_11415.LUT_INIT = 16'he4aa;
    SB_DFF i272_273 (.Q(\REG.mem_2_14 ), .C(FIFO_CLK_c), .D(n4959));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4076_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_33_1 ), .O(n5459));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4076_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i35_2_lut_3_lut (.I0(n11), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n35));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i35_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i4107_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_34_15 ), .O(n5490));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4107_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i269_270 (.Q(\REG.mem_2_13 ), .C(FIFO_CLK_c), .D(n4958));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4075_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_33_0 ), .O(n5458));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4075_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12779_bdd_4_lut (.I0(n12779), .I1(\REG.mem_45_12 ), .I2(\REG.mem_44_12 ), 
            .I3(rd_addr_r_c[1]), .O(n12782));
    defparam n12779_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i266_267 (.Q(\REG.mem_2_12 ), .C(FIFO_CLK_c), .D(n4957));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13433_bdd_4_lut (.I0(n13433), .I1(n11445), .I2(n11444), .I3(rd_addr_r_c[2]), 
            .O(n11583));
    defparam n13433_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i82_2_lut_3_lut_4_lut (.I0(n17_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n59));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i82_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_DFF i263_264 (.Q(\REG.mem_2_11 ), .C(FIFO_CLK_c), .D(n4956));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wr_addr_r_6__I_0_141_7_lut (.I0(GND_net), .I1(wr_addr_r[5]), 
            .I2(GND_net), .I3(n10137), .O(wr_addr_p1_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF i260_261 (.Q(\REG.mem_2_10 ), .C(FIFO_CLK_c), .D(n4955));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i81_2_lut_3_lut_4_lut (.I0(n17_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n27));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i81_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i4106_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_34_14 ), .O(n5489));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4106_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4436_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_53_15 ), .O(n5819));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4436_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4105_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_34_13 ), .O(n5488));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4105_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4435_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_53_14 ), .O(n5818));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4435_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4434_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_53_13 ), .O(n5817));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4434_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4433_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_53_12 ), .O(n5816));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4433_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4104_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_34_12 ), .O(n5487));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4104_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4432_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_53_11 ), .O(n5815));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4432_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4431_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_53_10 ), .O(n5814));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4431_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4103_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_34_11 ), .O(n5486));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4103_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11400 (.I0(rd_addr_r_c[1]), .I1(n11537), 
            .I2(n11538), .I3(rd_addr_r_c[2]), .O(n13427));
    defparam rd_addr_r_1__bdd_4_lut_11400.LUT_INIT = 16'he4aa;
    SB_LUT4 i4430_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_53_9 ), .O(n5813));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4430_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4429_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_53_8 ), .O(n5812));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4429_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i257_258 (.Q(\REG.mem_2_9 ), .C(FIFO_CLK_c), .D(n4954));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4102_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_34_10 ), .O(n5485));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4102_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9684_3_lut (.I0(\REG.mem_32_1 ), .I1(\REG.mem_33_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11522));
    defparam i9684_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i254_255 (.Q(\REG.mem_2_8 ), .C(FIFO_CLK_c), .D(n4953));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i17_2_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n17_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i17_2_lut.LUT_INIT = 16'h8888;
    SB_DFF i251_252 (.Q(\REG.mem_2_7 ), .C(FIFO_CLK_c), .D(n4952));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13427_bdd_4_lut (.I0(n13427), .I1(n11535), .I2(n11534), .I3(rd_addr_r_c[2]), 
            .O(n11586));
    defparam n13427_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i248_249 (.Q(\REG.mem_2_6 ), .C(FIFO_CLK_c), .D(n4951));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4428_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_53_7 ), .O(n5811));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4428_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4101_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_34_9 ), .O(n5484));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4101_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4100_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_34_8 ), .O(n5483));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4100_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11395 (.I0(rd_addr_r_c[1]), .I1(n11546), 
            .I2(n11547), .I3(rd_addr_r_c[2]), .O(n13421));
    defparam rd_addr_r_1__bdd_4_lut_11395.LUT_INIT = 16'he4aa;
    SB_LUT4 i9685_3_lut (.I0(\REG.mem_34_1 ), .I1(\REG.mem_35_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11523));
    defparam i9685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4427_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_53_6 ), .O(n5810));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4427_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4099_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_34_7 ), .O(n5482));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4099_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9574_3_lut (.I0(\REG.mem_34_7 ), .I1(\REG.mem_35_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11412));
    defparam i9574_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9573_3_lut (.I0(\REG.mem_32_7 ), .I1(\REG.mem_33_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11411));
    defparam i9573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9447_3_lut (.I0(\REG.mem_4_0 ), .I1(\REG.mem_5_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11285));
    defparam i9447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9448_3_lut (.I0(\REG.mem_6_0 ), .I1(\REG.mem_7_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11286));
    defparam i9448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4426_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_53_5 ), .O(n5809));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4426_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9445_3_lut (.I0(\REG.mem_2_0 ), .I1(\REG.mem_3_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11283));
    defparam i9445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9444_3_lut (.I0(\REG.mem_0_0 ), .I1(\REG.mem_1_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11282));
    defparam i9444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9651_3_lut (.I0(\REG.mem_36_10 ), .I1(\REG.mem_37_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11489));
    defparam i9651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9652_3_lut (.I0(\REG.mem_38_10 ), .I1(\REG.mem_39_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11490));
    defparam i9652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4425_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_53_4 ), .O(n5808));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4425_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9640_3_lut (.I0(\REG.mem_34_10 ), .I1(\REG.mem_35_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11478));
    defparam i9640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9639_3_lut (.I0(\REG.mem_32_10 ), .I1(\REG.mem_33_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11477));
    defparam i9639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9612_3_lut (.I0(\REG.mem_20_10 ), .I1(\REG.mem_21_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11450));
    defparam i9612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9613_3_lut (.I0(\REG.mem_22_10 ), .I1(\REG.mem_23_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11451));
    defparam i9613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4424_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_53_3 ), .O(n5807));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4424_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9610_3_lut (.I0(\REG.mem_18_10 ), .I1(\REG.mem_19_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11448));
    defparam i9610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9609_3_lut (.I0(\REG.mem_16_10 ), .I1(\REG.mem_17_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11447));
    defparam i9609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9405_3_lut (.I0(\REG.mem_4_7 ), .I1(\REG.mem_5_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11243));
    defparam i9405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9406_3_lut (.I0(\REG.mem_6_7 ), .I1(\REG.mem_7_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11244));
    defparam i9406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10083_3_lut (.I0(n12710), .I1(n12632), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11921));
    defparam i10083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10084_3_lut (.I0(n12512), .I1(n12410), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11922));
    defparam i10084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10063_3_lut (.I0(n12920), .I1(n12782), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11901));
    defparam i10063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10062_3_lut (.I0(n13004), .I1(n12974), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11900));
    defparam i10062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4423_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_53_2 ), .O(n5806));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4423_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9364_3_lut (.I0(\REG.mem_2_7 ), .I1(\REG.mem_3_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11202));
    defparam i9364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9363_3_lut (.I0(\REG.mem_0_7 ), .I1(\REG.mem_1_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11201));
    defparam i9363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4422_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_53_1 ), .O(n5805));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4422_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9585_3_lut (.I0(\REG.mem_4_10 ), .I1(\REG.mem_5_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11423));
    defparam i9585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9586_3_lut (.I0(\REG.mem_6_10 ), .I1(\REG.mem_7_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11424));
    defparam i9586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9577_3_lut (.I0(\REG.mem_2_10 ), .I1(\REG.mem_3_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11415));
    defparam i9577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9576_3_lut (.I0(\REG.mem_0_10 ), .I1(\REG.mem_1_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11414));
    defparam i9576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4421_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_53_0 ), .O(n5804));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4421_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9634_3_lut (.I0(n13388), .I1(n13202), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11472));
    defparam i9634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9622_3_lut (.I0(n13472), .I1(n12776), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11460));
    defparam i9622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9564_3_lut (.I0(\REG.mem_52_5 ), .I1(\REG.mem_53_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11402));
    defparam i9564_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9565_3_lut (.I0(\REG.mem_54_5 ), .I1(\REG.mem_55_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11403));
    defparam i9565_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9547_3_lut (.I0(\REG.mem_50_5 ), .I1(\REG.mem_51_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11385));
    defparam i9547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9546_3_lut (.I0(\REG.mem_48_5 ), .I1(\REG.mem_49_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11384));
    defparam i9546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i80_2_lut_3_lut_4_lut (.I0(n15_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n60));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i80_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i79_2_lut_3_lut_4_lut (.I0(n15_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n28));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i79_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i3_2_lut (.I0(\rd_addr_nxt_c_6__N_498[2] ), 
            .I1(\rd_addr_nxt_c_6__N_498[3] ), .I2(GND_net), .I3(GND_net), 
            .O(rd_grey_w[2]));   // src/fifo_dc_32_lut_gen.v(504[28:66])
    defparam rd_addr_nxt_c_6__I_0_152_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4420_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_52_15 ), .O(n5803));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4420_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10067_3_lut (.I0(n13424), .I1(n11904), .I2(rd_addr_r_c[3]), 
            .I3(GND_net), .O(n11905));
    defparam i10067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10066_3_lut (.I0(n13442), .I1(n13358), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11904));
    defparam i10066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4419_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_52_14 ), .O(n5802));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4419_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9366_3_lut (.I0(\REG.mem_20_5 ), .I1(\REG.mem_21_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11204));
    defparam i9366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9367_3_lut (.I0(\REG.mem_22_5 ), .I1(\REG.mem_23_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11205));
    defparam i9367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9325_3_lut (.I0(\REG.mem_18_5 ), .I1(\REG.mem_19_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11163));
    defparam i9325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9324_3_lut (.I0(\REG.mem_16_5 ), .I1(\REG.mem_17_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11162));
    defparam i9324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4418_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_52_13 ), .O(n5801));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4418_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4417_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_52_12 ), .O(n5800));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4417_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4416_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_52_11 ), .O(n5799));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4416_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9234_3_lut (.I0(\REG.mem_4_5 ), .I1(\REG.mem_5_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11072));
    defparam i9234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9235_3_lut (.I0(\REG.mem_6_5 ), .I1(\REG.mem_7_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11073));
    defparam i9235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4415_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_52_10 ), .O(n5798));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4415_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i47_2_lut_3_lut_4_lut (.I0(n12_adj_33), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n47_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i47_2_lut_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 EnabledDecoder_2_i49_2_lut_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n49_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i49_2_lut_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i4414_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_52_9 ), .O(n5797));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4414_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10098_3_lut (.I0(\REG.mem_60_8 ), .I1(\REG.mem_61_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11936));
    defparam i10098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10099_3_lut (.I0(\REG.mem_62_8 ), .I1(\REG.mem_63_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11937));
    defparam i10099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9199_3_lut (.I0(\REG.mem_2_5 ), .I1(\REG.mem_3_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11037));
    defparam i9199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9198_3_lut (.I0(\REG.mem_0_5 ), .I1(\REG.mem_1_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11036));
    defparam i9198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10036_3_lut (.I0(\REG.mem_58_8 ), .I1(\REG.mem_59_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11874));
    defparam i10036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10035_3_lut (.I0(\REG.mem_56_8 ), .I1(\REG.mem_57_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11873));
    defparam i10035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_5__I_0_i6_2_lut_3_lut (.I0(wr_addr_r[5]), .I1(rp_sync2_r[5]), 
            .I2(rp_sync2_r[6]), .I3(GND_net), .O(n6_adj_37));   // src/fifo_dc_32_lut_gen.v(295[31:67])
    defparam wr_addr_r_5__I_0_i6_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4413_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_52_8 ), .O(n5796));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4413_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut (.I0(rp_sync2_r[2]), .I1(rp_sync2_r[3]), .I2(rp_sync_w[4]), 
            .I3(GND_net), .O(rp_sync_w[2]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_39 (.I0(rp_sync2_r[0]), .I1(rp_sync2_r[1]), 
            .I2(rp_sync_w[2]), .I3(GND_net), .O(rp_sync_w[0]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_3_lut_adj_39.LUT_INIT = 16'h9696;
    SB_LUT4 i4098_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_34_6 ), .O(n5481));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4098_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_fifo_en_w_I_0_158_2_lut_3_lut (.I0(DEBUG_3_c), .I1(get_next_word), 
            .I2(\genblk16.rd_prev_r ), .I3(GND_net), .O(t_rd_fifo_en_w));   // src/fifo_dc_32_lut_gen.v(747[41:67])
    defparam rd_fifo_en_w_I_0_158_2_lut_3_lut.LUT_INIT = 16'hf4f4;
    SB_LUT4 i10089_3_lut (.I0(\REG.mem_60_15 ), .I1(\REG.mem_61_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11927));
    defparam i10089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10090_3_lut (.I0(\REG.mem_62_15 ), .I1(\REG.mem_63_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11928));
    defparam i10090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10081_3_lut (.I0(\REG.mem_58_15 ), .I1(\REG.mem_59_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11919));
    defparam i10081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10080_3_lut (.I0(\REG.mem_56_15 ), .I1(\REG.mem_57_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11918));
    defparam i10080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4097_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_34_5 ), .O(n5480));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4097_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4096_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_34_4 ), .O(n5479));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4096_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4412_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_52_7 ), .O(n5795));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4412_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4411_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_52_6 ), .O(n5794));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4411_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4410_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_52_5 ), .O(n5793));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4410_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4409_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_52_4 ), .O(n5792));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4409_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i57_2_lut_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n57_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i57_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i9441_3_lut (.I0(\REG.mem_36_9 ), .I1(\REG.mem_37_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11279));
    defparam i9441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9442_3_lut (.I0(\REG.mem_38_9 ), .I1(\REG.mem_39_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11280));
    defparam i9442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9415_3_lut (.I0(\REG.mem_34_9 ), .I1(\REG.mem_35_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11253));
    defparam i9415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9414_3_lut (.I0(\REG.mem_32_9 ), .I1(\REG.mem_33_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11252));
    defparam i9414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9372_3_lut (.I0(\REG.mem_20_9 ), .I1(\REG.mem_21_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11210));
    defparam i9372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9373_3_lut (.I0(\REG.mem_22_9 ), .I1(\REG.mem_23_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11211));
    defparam i9373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9349_3_lut (.I0(\REG.mem_18_9 ), .I1(\REG.mem_19_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11187));
    defparam i9349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9348_3_lut (.I0(\REG.mem_16_9 ), .I1(\REG.mem_17_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11186));
    defparam i9348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i59_2_lut_3_lut_4_lut (.I0(n11), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n59_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i59_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i9_2_lut_3_lut_4_lut (.I0(DEBUG_5_c), .I1(full_o), 
            .I2(wr_addr_r[0]), .I3(wr_addr_r[1]), .O(n9));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i9_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i4408_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_52_3 ), .O(n5791));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4408_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i42_2_lut_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n42_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i42_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i4095_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_34_3 ), .O(n5478));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4095_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4407_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_52_2 ), .O(n5790));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4407_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9051_4_lut_4_lut (.I0(rd_addr_r_c[1]), .I1(rd_addr_r_c[2]), 
            .I2(wp_sync2_r[1]), .I3(wp_sync_w[2]), .O(n10887));
    defparam i9051_4_lut_4_lut.LUT_INIT = 16'hb7de;
    SB_LUT4 i1_2_lut_3_lut_adj_40 (.I0(wp_sync2_r[4]), .I1(wp_sync2_r[6]), 
            .I2(wp_sync2_r[5]), .I3(GND_net), .O(wp_sync_w[4]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_adj_40.LUT_INIT = 16'h9696;
    SB_LUT4 i9594_3_lut (.I0(\REG.mem_60_5 ), .I1(\REG.mem_61_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11432));
    defparam i9594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9595_3_lut (.I0(\REG.mem_62_5 ), .I1(\REG.mem_63_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11433));
    defparam i9595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_41 (.I0(wp_sync2_r[0]), .I1(wp_sync2_r[1]), 
            .I2(wp_sync_w[2]), .I3(GND_net), .O(wp_sync_w[0]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_adj_41.LUT_INIT = 16'h9696;
    SB_LUT4 EnabledDecoder_2_i63_2_lut_3_lut_4_lut (.I0(n12_adj_33), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n63));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i63_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_3_lut_adj_42 (.I0(wp_sync2_r[2]), .I1(wp_sync2_r[3]), 
            .I2(wp_sync_w[4]), .I3(GND_net), .O(wp_sync_w[2]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_adj_42.LUT_INIT = 16'h9696;
    SB_LUT4 i9583_3_lut (.I0(\REG.mem_58_5 ), .I1(\REG.mem_59_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11421));
    defparam i9583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9582_3_lut (.I0(\REG.mem_56_5 ), .I1(\REG.mem_57_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11420));
    defparam i9582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4406_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_52_1 ), .O(n5789));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4406_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i65_2_lut_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n65));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i65_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i9655_3_lut (.I0(n12464), .I1(n12344), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11493));
    defparam i9655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9654_3_lut (.I0(n12890), .I1(n12584), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11492));
    defparam i9654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4405_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_52_0 ), .O(n5788));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4405_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9737_3_lut (.I0(n13058), .I1(n11574), .I2(rd_addr_r_c[3]), 
            .I3(GND_net), .O(n11575));
    defparam i9737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9736_3_lut (.I0(n12998), .I1(n12926), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11574));
    defparam i9736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10076_3_lut (.I0(n13454), .I1(n11913), .I2(rd_addr_r_c[3]), 
            .I3(GND_net), .O(n11914));
    defparam i10076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10075_3_lut (.I0(n13784), .I1(n13256), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11913));
    defparam i10075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9411_3_lut (.I0(n12302), .I1(n13664), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11249));
    defparam i9411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9396_3_lut (.I0(\REG.mem_52_4 ), .I1(\REG.mem_53_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11234));
    defparam i9396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9397_3_lut (.I0(\REG.mem_54_4 ), .I1(\REG.mem_55_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11235));
    defparam i9397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9388_3_lut (.I0(\REG.mem_50_4 ), .I1(\REG.mem_51_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11226));
    defparam i9388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9387_3_lut (.I0(\REG.mem_48_4 ), .I1(\REG.mem_49_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11225));
    defparam i9387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9375_3_lut (.I0(\REG.mem_36_4 ), .I1(\REG.mem_37_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11213));
    defparam i9375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9376_3_lut (.I0(\REG.mem_38_4 ), .I1(\REG.mem_39_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11214));
    defparam i9376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9370_3_lut (.I0(\REG.mem_34_4 ), .I1(\REG.mem_35_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11208));
    defparam i9370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9369_3_lut (.I0(\REG.mem_32_4 ), .I1(\REG.mem_33_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11207));
    defparam i9369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9351_3_lut (.I0(\REG.mem_20_4 ), .I1(\REG.mem_21_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11189));
    defparam i9351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9352_3_lut (.I0(\REG.mem_22_4 ), .I1(\REG.mem_23_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11190));
    defparam i9352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9340_3_lut (.I0(\REG.mem_18_4 ), .I1(\REG.mem_19_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11178));
    defparam i9340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9339_3_lut (.I0(\REG.mem_16_4 ), .I1(\REG.mem_17_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11177));
    defparam i9339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9190_3_lut (.I0(n12392), .I1(n12356), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11028));
    defparam i9190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9189_3_lut (.I0(n12626), .I1(n12530), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11027));
    defparam i9189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9597_3_lut (.I0(\REG.mem_12_10 ), .I1(\REG.mem_13_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11435));
    defparam i9597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9598_3_lut (.I0(\REG.mem_14_10 ), .I1(\REG.mem_15_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11436));
    defparam i9598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9589_3_lut (.I0(\REG.mem_10_10 ), .I1(\REG.mem_11_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11427));
    defparam i9589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9588_3_lut (.I0(\REG.mem_8_10 ), .I1(\REG.mem_9_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11426));
    defparam i9588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i45_2_lut_3_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n45));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i45_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i78_2_lut_3_lut_4_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n61));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i78_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i77_2_lut_3_lut_4_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n29));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i77_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i4404_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_51_15 ), .O(n5787));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4404_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4403_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_51_14 ), .O(n5786));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4403_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4402_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_51_13 ), .O(n5785));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4402_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4401_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_51_12 ), .O(n5784));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4401_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4400_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_51_11 ), .O(n5783));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4400_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9630_3_lut (.I0(\REG.mem_28_10 ), .I1(\REG.mem_29_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11468));
    defparam i9630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9631_3_lut (.I0(\REG.mem_30_10 ), .I1(\REG.mem_31_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11469));
    defparam i9631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4399_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_51_10 ), .O(n5782));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4399_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4398_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_51_9 ), .O(n5781));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4398_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4397_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_51_8 ), .O(n5780));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4397_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4396_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_51_7 ), .O(n5779));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4396_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9619_3_lut (.I0(\REG.mem_26_10 ), .I1(\REG.mem_27_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11457));
    defparam i9619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9618_3_lut (.I0(\REG.mem_24_10 ), .I1(\REG.mem_25_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11456));
    defparam i9618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9669_3_lut (.I0(\REG.mem_44_10 ), .I1(\REG.mem_45_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11507));
    defparam i9669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9670_3_lut (.I0(\REG.mem_46_10 ), .I1(\REG.mem_47_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11508));
    defparam i9670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9658_3_lut (.I0(\REG.mem_42_10 ), .I1(\REG.mem_43_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11496));
    defparam i9658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9657_3_lut (.I0(\REG.mem_40_10 ), .I1(\REG.mem_41_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11495));
    defparam i9657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10050_3_lut (.I0(n13322), .I1(n13262), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11888));
    defparam i10050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10051_3_lut (.I0(n13196), .I1(n13130), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11889));
    defparam i10051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10039_3_lut (.I0(n13460), .I1(n13382), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11877));
    defparam i10039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10077_3_lut (.I0(\REG.mem_28_14 ), .I1(\REG.mem_29_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11915));
    defparam i10077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10078_3_lut (.I0(\REG.mem_30_14 ), .I1(\REG.mem_31_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11916));
    defparam i10078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10054_3_lut (.I0(\REG.mem_26_14 ), .I1(\REG.mem_27_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11892));
    defparam i10054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10053_3_lut (.I0(\REG.mem_24_14 ), .I1(\REG.mem_25_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11891));
    defparam i10053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10188_3_lut (.I0(\REG.mem_20_13 ), .I1(\REG.mem_21_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12026));
    defparam i10188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10189_3_lut (.I0(\REG.mem_22_13 ), .I1(\REG.mem_23_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12027));
    defparam i10189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10146_3_lut (.I0(\REG.mem_36_14 ), .I1(\REG.mem_37_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11984));
    defparam i10146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10147_3_lut (.I0(\REG.mem_38_14 ), .I1(\REG.mem_39_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11985));
    defparam i10147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10135_3_lut (.I0(\REG.mem_18_13 ), .I1(\REG.mem_19_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11973));
    defparam i10135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10134_3_lut (.I0(\REG.mem_16_13 ), .I1(\REG.mem_17_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11972));
    defparam i10134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10141_3_lut (.I0(\REG.mem_34_14 ), .I1(\REG.mem_35_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11979));
    defparam i10141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10140_3_lut (.I0(\REG.mem_32_14 ), .I1(\REG.mem_33_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11978));
    defparam i10140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10183_3_lut (.I0(n13622), .I1(n13448), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n12021));
    defparam i10183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10165_3_lut (.I0(n13604), .I1(n12704), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n12003));
    defparam i10165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10164_3_lut (.I0(n13490), .I1(n13658), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n12002));
    defparam i10164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9627_3_lut (.I0(\REG.mem_44_7 ), .I1(\REG.mem_45_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11465));
    defparam i9627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9628_3_lut (.I0(\REG.mem_46_7 ), .I1(\REG.mem_47_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11466));
    defparam i9628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9607_3_lut (.I0(\REG.mem_42_7 ), .I1(\REG.mem_43_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11445));
    defparam i9607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9606_3_lut (.I0(\REG.mem_40_7 ), .I1(\REG.mem_41_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11444));
    defparam i9606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i11_2_lut_3_lut_4_lut (.I0(DEBUG_5_c), .I1(full_o), 
            .I2(wr_addr_r[0]), .I3(wr_addr_r[1]), .O(n11));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i9699_3_lut (.I0(\REG.mem_60_10 ), .I1(\REG.mem_61_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11537));
    defparam i9699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9700_3_lut (.I0(\REG.mem_62_10 ), .I1(\REG.mem_63_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11538));
    defparam i9700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i12_2_lut_3_lut_4_lut (.I0(DEBUG_5_c), .I1(full_o), 
            .I2(wr_addr_r[0]), .I3(wr_addr_r[1]), .O(n12_adj_33));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i12_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i9697_3_lut (.I0(\REG.mem_58_10 ), .I1(\REG.mem_59_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11535));
    defparam i9697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9696_3_lut (.I0(\REG.mem_56_10 ), .I1(\REG.mem_57_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11534));
    defparam i9696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i43_2_lut_3_lut_4_lut (.I0(n11), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n43));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i43_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i9708_3_lut (.I0(\REG.mem_36_1 ), .I1(\REG.mem_37_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11546));
    defparam i9708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9709_3_lut (.I0(\REG.mem_38_1 ), .I1(\REG.mem_39_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11547));
    defparam i9709_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module clock
//

module clock (GND_net, VCC_net, ICE_SYSCLK_c, pll_clk_unbuf) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    input ICE_SYSCLK_c;
    output pll_clk_unbuf;
    
    
    SB_PLL40_CORE pll_config (.REFERENCECLK(ICE_SYSCLK_c), .PLLOUTGLOBAL(pll_clk_unbuf), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=222, LSE_RLINE=228 */ ;   // src/top.v(222[7] 228[3])
    defparam pll_config.FEEDBACK_PATH = "SIMPLE";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll_config.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll_config.FDA_FEEDBACK = 0;
    defparam pll_config.FDA_RELATIVE = 0;
    defparam pll_config.PLLOUT_SELECT = "GENCLK";
    defparam pll_config.DIVR = 4'b0001;
    defparam pll_config.DIVF = 7'b1010010;
    defparam pll_config.DIVQ = 3'b100;
    defparam pll_config.FILTER_RANGE = 3'b001;
    defparam pll_config.ENABLE_ICEGATE = 1'b0;
    defparam pll_config.TEST_MODE = 1'b0;
    defparam pll_config.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=20) 
//

module \uart_rx(CLKS_PER_BIT=20)  (r_SM_Main, SLM_CLK_c, r_Rx_Data, GND_net, 
            n4, n4_adj_1, n6105, pc_data_rx, n10406, VCC_net, debug_led3, 
            n7473, n6082, n6081, n6079, n6078, n6077, n6075, n6074, 
            \r_SM_Main_2__N_765[2] , n4_adj_2, n10345, UART_RX_c, n4248, 
            n4253) /* synthesis syn_module_defined=1 */ ;
    output [2:0]r_SM_Main;
    input SLM_CLK_c;
    output r_Rx_Data;
    input GND_net;
    output n4;
    output n4_adj_1;
    input n6105;
    output [7:0]pc_data_rx;
    input n10406;
    input VCC_net;
    output debug_led3;
    output n7473;
    input n6082;
    input n6081;
    input n6079;
    input n6078;
    input n6077;
    input n6075;
    input n6074;
    output \r_SM_Main_2__N_765[2] ;
    output n4_adj_2;
    output n10345;
    input UART_RX_c;
    output n4248;
    output n4253;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n3, r_Rx_Data_R;
    wire [9:0]n45;
    
    wire n6700;
    wire [9:0]r_Clock_Count;   // src/uart_rx.v(32[17:30])
    
    wire n6691, n151, n6072;
    wire [2:0]r_Bit_Index;   // src/uart_rx.v(33[17:28])
    
    wire n10448, n4367, n55_adj_18, n145, n3_adj_19, n10213, n10212, 
        n10211, n10210, n13, n125, n10209, n10208, n10207;
    wire [2:0]n340;
    
    wire n4676, n149, n10206, n4_adj_20, n140, n6, n8, n6725, 
        n6710, n10205;
    
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(SLM_CLK_c), .D(n3), .R(r_SM_Main[2]));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(SLM_CLK_c), .D(r_Rx_Data_R));   // src/uart_rx.v(41[10] 45[8])
    SB_DFFESR r_Clock_Count_1191__i0 (.Q(r_Clock_Count[0]), .C(SLM_CLK_c), 
            .E(n6700), .D(n45[0]), .R(n6691));   // src/uart_rx.v(120[34:51])
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(n151), .I2(GND_net), .I3(GND_net), 
            .O(n6072));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_140_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // src/uart_rx.v(97[17:39])
    defparam equal_140_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_137_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // src/uart_rx.v(97[17:39])
    defparam equal_137_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFF r_Rx_Byte_i0 (.Q(pc_data_rx[0]), .C(SLM_CLK_c), .D(n6105));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Rx_DV_52 (.Q(debug_led3), .C(SLM_CLK_c), .E(VCC_net), .D(n10406));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i6110_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n7473));
    defparam i6110_2_lut.LUT_INIT = 16'h8888;
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n10448));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(pc_data_rx[7]), .C(SLM_CLK_c), .D(n6082));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(pc_data_rx[6]), .C(SLM_CLK_c), .D(n6081));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(pc_data_rx[5]), .C(SLM_CLK_c), .D(n6079));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(pc_data_rx[4]), .C(SLM_CLK_c), .D(n6078));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(pc_data_rx[3]), .C(SLM_CLK_c), .D(n6077));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(pc_data_rx[2]), .C(SLM_CLK_c), .D(n6075));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(pc_data_rx[1]), .C(SLM_CLK_c), .D(n6074));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(SLM_CLK_c), .D(n6072));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_4_lut (.I0(\r_SM_Main_2__N_765[2] ), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main[2]), .O(n4367));
    defparam i2_4_lut.LUT_INIT = 16'h0023;
    SB_LUT4 i12_3_lut (.I0(n4367), .I1(r_Bit_Index[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n10448));   // src/uart_rx.v(36[17:26])
    defparam i12_3_lut.LUT_INIT = 16'h6464;
    SB_LUT4 equal_141_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // src/uart_rx.v(97[17:39])
    defparam equal_141_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[0]), .I1(n151), .I2(n4_adj_2), .I3(r_Bit_Index[0]), 
            .O(n10345));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(SLM_CLK_c), .D(UART_RX_c));   // src/uart_rx.v(41[10] 45[8])
    SB_LUT4 i1_2_lut_3_lut (.I0(r_SM_Main[0]), .I1(n151), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n4248));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_21 (.I0(r_SM_Main[0]), .I1(n151), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n4253));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_adj_21.LUT_INIT = 16'hbfbf;
    SB_LUT4 i1_2_lut_adj_22 (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_765[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n55_adj_18));
    defparam i1_2_lut_adj_22.LUT_INIT = 16'h8888;
    SB_LUT4 i5351_4_lut (.I0(r_Rx_Data), .I1(n55_adj_18), .I2(r_SM_Main[1]), 
            .I3(n145), .O(n3_adj_19));   // src/uart_rx.v(36[17:26])
    defparam i5351_4_lut.LUT_INIT = 16'h3530;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(SLM_CLK_c), .D(n3_adj_19), 
            .R(r_SM_Main[2]));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_Clock_Count_1191_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[9]), .I3(n10213), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1191_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n10212), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1191_add_4_10 (.CI(n10212), .I0(GND_net), .I1(r_Clock_Count[8]), 
            .CO(n10213));
    SB_DFFESR r_Clock_Count_1191__i9 (.Q(r_Clock_Count[9]), .C(SLM_CLK_c), 
            .E(n6700), .D(n45[9]), .R(n6691));   // src/uart_rx.v(120[34:51])
    SB_LUT4 r_Clock_Count_1191_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n10211), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1191_add_4_9 (.CI(n10211), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n10212));
    SB_DFFESR r_Clock_Count_1191__i8 (.Q(r_Clock_Count[8]), .C(SLM_CLK_c), 
            .E(n6700), .D(n45[8]), .R(n6691));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1191__i7 (.Q(r_Clock_Count[7]), .C(SLM_CLK_c), 
            .E(n6700), .D(n45[7]), .R(n6691));   // src/uart_rx.v(120[34:51])
    SB_LUT4 r_Clock_Count_1191_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n10210), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main[0]), .I2(n13), .I3(GND_net), 
            .O(n125));   // src/uart_rx.v(30[17:26])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i10396_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[2]), .I2(n145), 
            .I3(r_SM_Main[1]), .O(n6700));
    defparam i10396_4_lut.LUT_INIT = 16'h3313;
    SB_CARRY r_Clock_Count_1191_add_4_8 (.CI(n10210), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n10211));
    SB_LUT4 r_Clock_Count_1191_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n10209), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1191_add_4_7 (.CI(n10209), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n10210));
    SB_DFFESR r_Clock_Count_1191__i6 (.Q(r_Clock_Count[6]), .C(SLM_CLK_c), 
            .E(n6700), .D(n45[6]), .R(n6691));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1191__i5 (.Q(r_Clock_Count[5]), .C(SLM_CLK_c), 
            .E(n6700), .D(n45[5]), .R(n6691));   // src/uart_rx.v(120[34:51])
    SB_LUT4 r_Clock_Count_1191_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n10208), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1191_add_4_6 (.CI(n10208), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n10209));
    SB_DFFESR r_Clock_Count_1191__i4 (.Q(r_Clock_Count[4]), .C(SLM_CLK_c), 
            .E(n6700), .D(n45[4]), .R(n6691));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1191__i3 (.Q(r_Clock_Count[3]), .C(SLM_CLK_c), 
            .E(n6700), .D(n45[3]), .R(n6691));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1191__i2 (.Q(r_Clock_Count[2]), .C(SLM_CLK_c), 
            .E(n6700), .D(n45[2]), .R(n6691));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1191__i1 (.Q(r_Clock_Count[1]), .C(SLM_CLK_c), 
            .E(n6700), .D(n45[1]), .R(n6691));   // src/uart_rx.v(120[34:51])
    SB_LUT4 r_Clock_Count_1191_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n10207), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1191_add_4_5 (.CI(n10207), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n10208));
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(SLM_CLK_c), .E(n4367), 
            .D(n340[1]), .R(n4676));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1350_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n340[2]));   // src/uart_rx.v(49[10] 144[8])
    defparam i1350_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(n149));   // src/uart_rx.v(49[10] 144[8])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 r_Clock_Count_1191_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n10206), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_23 (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), 
            .I2(r_Clock_Count[1]), .I3(GND_net), .O(n4_adj_20));   // src/uart_rx.v(118[17:47])
    defparam i1_3_lut_adj_23.LUT_INIT = 16'hecec;
    SB_LUT4 i1_4_lut (.I0(r_Clock_Count[4]), .I1(n140), .I2(r_Clock_Count[3]), 
            .I3(n4_adj_20), .O(\r_SM_Main_2__N_765[2] ));   // src/uart_rx.v(32[17:30])
    defparam i1_4_lut.LUT_INIT = 16'heeec;
    SB_LUT4 i1_2_lut_adj_24 (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[7]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // src/uart_rx.v(32[17:30])
    defparam i1_2_lut_adj_24.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[6]), .I2(r_Clock_Count[9]), 
            .I3(n6), .O(n140));   // src/uart_rx.v(32[17:30])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_25 (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[1]), 
            .I2(r_Clock_Count[3]), .I3(r_Clock_Count[4]), .O(n8));
    defparam i3_4_lut_adj_25.LUT_INIT = 16'hffdf;
    SB_LUT4 i4_3_lut (.I0(n140), .I1(n8), .I2(r_Clock_Count[2]), .I3(GND_net), 
            .O(n13));
    defparam i4_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_26 (.I0(r_SM_Main[0]), .I1(n13), .I2(GND_net), 
            .I3(GND_net), .O(n145));   // src/uart_rx.v(36[17:26])
    defparam i1_2_lut_adj_26.LUT_INIT = 16'h2222;
    SB_LUT4 i5343_3_lut (.I0(n149), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_765[2] ), 
            .I3(GND_net), .O(n6725));   // src/uart_rx.v(36[17:26])
    defparam i5343_3_lut.LUT_INIT = 16'h2c2c;
    SB_LUT4 i5344_3_lut (.I0(n6710), .I1(n6725), .I2(r_SM_Main[1]), .I3(GND_net), 
            .O(n3));   // src/uart_rx.v(36[17:26])
    defparam i5344_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY r_Clock_Count_1191_add_4_4 (.CI(n10206), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n10207));
    SB_LUT4 i5309_4_lut_4_lut (.I0(\r_SM_Main_2__N_765[2] ), .I1(r_SM_Main[2]), 
            .I2(n125), .I3(r_SM_Main[1]), .O(n6691));   // src/uart_rx.v(49[10] 144[8])
    defparam i5309_4_lut_4_lut.LUT_INIT = 16'h2203;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(SLM_CLK_c), .E(n4367), 
            .D(n340[2]), .R(n4676));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_Clock_Count_1191_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n10205), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_27 (.I0(\r_SM_Main_2__N_765[2] ), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n151));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_adj_27.LUT_INIT = 16'h2020;
    SB_CARRY r_Clock_Count_1191_add_4_3 (.CI(n10205), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n10206));
    SB_LUT4 r_Clock_Count_1191_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1191_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n10205));
    SB_LUT4 i5328_4_lut_3_lut (.I0(r_SM_Main[0]), .I1(n13), .I2(r_Rx_Data), 
            .I3(GND_net), .O(n6710));   // src/uart_rx.v(30[17:26])
    defparam i5328_4_lut_3_lut.LUT_INIT = 16'h8d8d;
    SB_LUT4 i1343_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n340[1]));   // src/uart_rx.v(102[36:51])
    defparam i1343_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3293_3_lut (.I0(n4367), .I1(r_SM_Main[1]), .I2(n149), .I3(GND_net), 
            .O(n4676));   // src/uart_rx.v(49[10] 144[8])
    defparam i3293_3_lut.LUT_INIT = 16'ha2a2;
    
endmodule
//
// Verilog Description of module FIFO_Quad_Word
//

module FIFO_Quad_Word (rd_fifo_en_w, \mem_LUT.data_raw_r[7] , SLM_CLK_c, 
            \mem_LUT.data_raw_r[6] , \mem_LUT.data_raw_r[5] , \mem_LUT.data_raw_r[0] , 
            \mem_LUT.data_raw_r[4] , \mem_LUT.data_raw_r[3] , rd_addr_r, 
            reset_all_w, n8, wr_addr_r, \mem_LUT.data_raw_r[2] , \mem_LUT.data_raw_r[1] , 
            GND_net, \rd_addr_p1_w[2] , n14025, n6127, VCC_net, \fifo_temp_output[1] , 
            n10430, is_tx_fifo_full_flag, n6088, \fifo_temp_output[0] , 
            \wr_addr_p1_w[2] , n1, n10226, n5989, n5311, \fifo_temp_output[4] , 
            n5314, \fifo_temp_output[5] , rx_buf_byte, n5868, n4882, 
            \fifo_temp_output[2] , n4887, \fifo_temp_output[3] , n5536, 
            \fifo_temp_output[6] , n5539, \fifo_temp_output[7] , n10786, 
            is_fifo_empty_flag, n4919, n4922, fifo_write_cmd, wr_fifo_en_w, 
            n4878, rd_fifo_en_prev_r, fifo_read_cmd) /* synthesis syn_module_defined=1 */ ;
    output rd_fifo_en_w;
    output \mem_LUT.data_raw_r[7] ;
    input SLM_CLK_c;
    output \mem_LUT.data_raw_r[6] ;
    output \mem_LUT.data_raw_r[5] ;
    output \mem_LUT.data_raw_r[0] ;
    output \mem_LUT.data_raw_r[4] ;
    output \mem_LUT.data_raw_r[3] ;
    output [2:0]rd_addr_r;
    input reset_all_w;
    input n8;
    output [2:0]wr_addr_r;
    output \mem_LUT.data_raw_r[2] ;
    output \mem_LUT.data_raw_r[1] ;
    input GND_net;
    output \rd_addr_p1_w[2] ;
    output n14025;
    input n6127;
    input VCC_net;
    output \fifo_temp_output[1] ;
    input n10430;
    output is_tx_fifo_full_flag;
    input n6088;
    output \fifo_temp_output[0] ;
    output \wr_addr_p1_w[2] ;
    output n1;
    output n10226;
    input n5989;
    input n5311;
    output \fifo_temp_output[4] ;
    input n5314;
    output \fifo_temp_output[5] ;
    input [7:0]rx_buf_byte;
    input n5868;
    input n4882;
    output \fifo_temp_output[2] ;
    input n4887;
    output \fifo_temp_output[3] ;
    input n5536;
    output \fifo_temp_output[6] ;
    input n5539;
    output \fifo_temp_output[7] ;
    input n10786;
    output is_fifo_empty_flag;
    input n4919;
    input n4922;
    input fifo_write_cmd;
    output wr_fifo_en_w;
    input n4878;
    output rd_fifo_en_prev_r;
    input fifo_read_cmd;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_2 lscc_fifo_inst (.rd_fifo_en_w(rd_fifo_en_w), 
            .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r[7] ), .SLM_CLK_c(SLM_CLK_c), 
            .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r[6] ), .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r[5] ), 
            .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r[0] ), .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r[4] ), 
            .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r[3] ), .rd_addr_r({rd_addr_r}), 
            .reset_all_w(reset_all_w), .n8(n8), .wr_addr_r({wr_addr_r}), 
            .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r[2] ), .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r[1] ), 
            .GND_net(GND_net), .\rd_addr_p1_w[2] (\rd_addr_p1_w[2] ), .n14025(n14025), 
            .n6127(n6127), .VCC_net(VCC_net), .\fifo_temp_output[1] (\fifo_temp_output[1] ), 
            .n10430(n10430), .is_tx_fifo_full_flag(is_tx_fifo_full_flag), 
            .n6088(n6088), .\fifo_temp_output[0] (\fifo_temp_output[0] ), 
            .\wr_addr_p1_w[2] (\wr_addr_p1_w[2] ), .n1(n1), .n10226(n10226), 
            .n5989(n5989), .n5311(n5311), .\fifo_temp_output[4] (\fifo_temp_output[4] ), 
            .n5314(n5314), .\fifo_temp_output[5] (\fifo_temp_output[5] ), 
            .rx_buf_byte({rx_buf_byte}), .n5868(n5868), .n4882(n4882), 
            .\fifo_temp_output[2] (\fifo_temp_output[2] ), .n4887(n4887), 
            .\fifo_temp_output[3] (\fifo_temp_output[3] ), .n5536(n5536), 
            .\fifo_temp_output[6] (\fifo_temp_output[6] ), .n5539(n5539), 
            .\fifo_temp_output[7] (\fifo_temp_output[7] ), .n10786(n10786), 
            .is_fifo_empty_flag(is_fifo_empty_flag), .n4919(n4919), .n4922(n4922), 
            .fifo_write_cmd(fifo_write_cmd), .wr_fifo_en_w(wr_fifo_en_w), 
            .n4878(n4878), .rd_fifo_en_prev_r(rd_fifo_en_prev_r), .fifo_read_cmd(fifo_read_cmd)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_quad_word_mod.v(20[37:380])
    
endmodule
//
// Verilog Description of module FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_2
//

module FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_2 (rd_fifo_en_w, 
            \mem_LUT.data_raw_r[7] , SLM_CLK_c, \mem_LUT.data_raw_r[6] , 
            \mem_LUT.data_raw_r[5] , \mem_LUT.data_raw_r[0] , \mem_LUT.data_raw_r[4] , 
            \mem_LUT.data_raw_r[3] , rd_addr_r, reset_all_w, n8, wr_addr_r, 
            \mem_LUT.data_raw_r[2] , \mem_LUT.data_raw_r[1] , GND_net, 
            \rd_addr_p1_w[2] , n14025, n6127, VCC_net, \fifo_temp_output[1] , 
            n10430, is_tx_fifo_full_flag, n6088, \fifo_temp_output[0] , 
            \wr_addr_p1_w[2] , n1, n10226, n5989, n5311, \fifo_temp_output[4] , 
            n5314, \fifo_temp_output[5] , rx_buf_byte, n5868, n4882, 
            \fifo_temp_output[2] , n4887, \fifo_temp_output[3] , n5536, 
            \fifo_temp_output[6] , n5539, \fifo_temp_output[7] , n10786, 
            is_fifo_empty_flag, n4919, n4922, fifo_write_cmd, wr_fifo_en_w, 
            n4878, rd_fifo_en_prev_r, fifo_read_cmd) /* synthesis syn_module_defined=1 */ ;
    output rd_fifo_en_w;
    output \mem_LUT.data_raw_r[7] ;
    input SLM_CLK_c;
    output \mem_LUT.data_raw_r[6] ;
    output \mem_LUT.data_raw_r[5] ;
    output \mem_LUT.data_raw_r[0] ;
    output \mem_LUT.data_raw_r[4] ;
    output \mem_LUT.data_raw_r[3] ;
    output [2:0]rd_addr_r;
    input reset_all_w;
    input n8;
    output [2:0]wr_addr_r;
    output \mem_LUT.data_raw_r[2] ;
    output \mem_LUT.data_raw_r[1] ;
    input GND_net;
    output \rd_addr_p1_w[2] ;
    output n14025;
    input n6127;
    input VCC_net;
    output \fifo_temp_output[1] ;
    input n10430;
    output is_tx_fifo_full_flag;
    input n6088;
    output \fifo_temp_output[0] ;
    output \wr_addr_p1_w[2] ;
    output n1;
    output n10226;
    input n5989;
    input n5311;
    output \fifo_temp_output[4] ;
    input n5314;
    output \fifo_temp_output[5] ;
    input [7:0]rx_buf_byte;
    input n5868;
    input n4882;
    output \fifo_temp_output[2] ;
    input n4887;
    output \fifo_temp_output[3] ;
    input n5536;
    output \fifo_temp_output[6] ;
    input n5539;
    output \fifo_temp_output[7] ;
    input n10786;
    output is_fifo_empty_flag;
    input n4919;
    input n4922;
    input fifo_write_cmd;
    output wr_fifo_en_w;
    input n4878;
    output rd_fifo_en_prev_r;
    input fifo_read_cmd;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [31:0]\mem_LUT.data_raw_r_31__N_1084 ;
    wire [2:0]n12;
    
    wire n2, \mem_LUT.mem_2_7 , \mem_LUT.mem_3_7 , n12587, \mem_LUT.mem_1_7 , 
        \mem_LUT.mem_0_7 , \mem_LUT.mem_2_6 , \mem_LUT.mem_3_6 , n12569, 
        \mem_LUT.mem_1_6 , \mem_LUT.mem_0_6 , \mem_LUT.mem_2_5 , \mem_LUT.mem_3_5 , 
        n12563, n6068, n6067, n6066, n6065, \mem_LUT.mem_3_4 , n6064, 
        \mem_LUT.mem_3_3 , n6063, \mem_LUT.mem_3_2 , n6062, \mem_LUT.mem_3_1 , 
        n6061, \mem_LUT.mem_3_0 , \mem_LUT.mem_1_5 , \mem_LUT.mem_0_5 , 
        \mem_LUT.mem_2_4 , n12557, n6053, n6052, n6051, n6050, n6049, 
        \mem_LUT.mem_2_3 , n6048, \mem_LUT.mem_2_2 , n6047, \mem_LUT.mem_2_1 , 
        n6046, \mem_LUT.mem_2_0 , n6040, n6039, n6038, n6037, \mem_LUT.mem_1_4 , 
        n6036, \mem_LUT.mem_1_3 , n6035, \mem_LUT.mem_1_2 , n6034, 
        \mem_LUT.mem_1_1 , \mem_LUT.mem_0_4 , n6033, \mem_LUT.mem_1_0 , 
        n6032, n6031, n6030, n6029, n6028, \mem_LUT.mem_0_3 , n6027, 
        \mem_LUT.mem_0_2 , n6026, \mem_LUT.mem_0_1 , n6025, \mem_LUT.mem_0_0 , 
        n12491, n3, n12485, n12473, n12437, n4;
    
    SB_DFFE \mem_LUT.data_raw_r__i8  (.Q(\mem_LUT.data_raw_r[7] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1084 [7]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i7  (.Q(\mem_LUT.data_raw_r[6] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1084 [6]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i6  (.Q(\mem_LUT.data_raw_r[5] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1084 [5]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i1  (.Q(\mem_LUT.data_raw_r[0] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1084 [0]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i5  (.Q(\mem_LUT.data_raw_r[4] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1084 [4]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i4  (.Q(\mem_LUT.data_raw_r[3] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1084 [3]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFSR rd_addr_r__i0 (.Q(rd_addr_r[0]), .C(SLM_CLK_c), .D(n12[0]), 
            .R(reset_all_w));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFSR wr_addr_r__i0 (.Q(wr_addr_r[0]), .C(SLM_CLK_c), .D(n8), .R(reset_all_w));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFE \mem_LUT.data_raw_r__i3  (.Q(\mem_LUT.data_raw_r[2] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1084 [2]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i2  (.Q(\mem_LUT.data_raw_r[1] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1084 [1]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_LUT4 wr_addr_p1_w_1__I_0_i2_2_lut_3_lut (.I0(wr_addr_r[1]), .I1(wr_addr_r[0]), 
            .I2(rd_addr_r[1]), .I3(GND_net), .O(n2));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam wr_addr_p1_w_1__I_0_i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1416_3_lut (.I0(rd_addr_r[2]), .I1(rd_addr_r[1]), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(\rd_addr_p1_w[2] ));   // src/fifo_quad_word_mod.v(71[47:65])
    defparam i1416_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1409_rep_150_2_lut (.I0(rd_addr_r[1]), .I1(rd_addr_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n14025));   // src/fifo_quad_word_mod.v(71[47:65])
    defparam i1409_rep_150_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 rd_addr_r_0__bdd_4_lut (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_7 ), 
            .I2(\mem_LUT.mem_3_7 ), .I3(rd_addr_r[1]), .O(n12587));
    defparam rd_addr_r_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n12587_bdd_4_lut (.I0(n12587), .I1(\mem_LUT.mem_1_7 ), .I2(\mem_LUT.mem_0_7 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1084 [7]));
    defparam n12587_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \mem_LUT.data_buff_r__i1  (.Q(\fifo_temp_output[1] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n6127));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE full_r_84 (.Q(is_tx_fifo_full_flag), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n10430));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFE \mem_LUT.data_buff_r__i0  (.Q(\fifo_temp_output[0] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n6088));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10697 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_6 ), 
            .I2(\mem_LUT.mem_3_6 ), .I3(rd_addr_r[1]), .O(n12569));
    defparam rd_addr_r_0__bdd_4_lut_10697.LUT_INIT = 16'he4aa;
    SB_LUT4 n12569_bdd_4_lut (.I0(n12569), .I1(\mem_LUT.mem_1_6 ), .I2(\mem_LUT.mem_0_6 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1084 [6]));
    defparam n12569_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10682 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_5 ), 
            .I2(\mem_LUT.mem_3_5 ), .I3(rd_addr_r[1]), .O(n12563));
    defparam rd_addr_r_0__bdd_4_lut_10682.LUT_INIT = 16'he4aa;
    SB_DFF i347_348 (.Q(\mem_LUT.mem_3_7 ), .C(SLM_CLK_c), .D(n6068));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i344_345 (.Q(\mem_LUT.mem_3_6 ), .C(SLM_CLK_c), .D(n6067));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i341_342 (.Q(\mem_LUT.mem_3_5 ), .C(SLM_CLK_c), .D(n6066));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i338_339 (.Q(\mem_LUT.mem_3_4 ), .C(SLM_CLK_c), .D(n6065));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i335_336 (.Q(\mem_LUT.mem_3_3 ), .C(SLM_CLK_c), .D(n6064));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i332_333 (.Q(\mem_LUT.mem_3_2 ), .C(SLM_CLK_c), .D(n6063));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i329_330 (.Q(\mem_LUT.mem_3_1 ), .C(SLM_CLK_c), .D(n6062));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i326_327 (.Q(\mem_LUT.mem_3_0 ), .C(SLM_CLK_c), .D(n6061));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 n12563_bdd_4_lut (.I0(n12563), .I1(\mem_LUT.mem_1_5 ), .I2(\mem_LUT.mem_0_5 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1084 [5]));
    defparam n12563_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10677 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_4 ), 
            .I2(\mem_LUT.mem_3_4 ), .I3(rd_addr_r[1]), .O(n12557));
    defparam rd_addr_r_0__bdd_4_lut_10677.LUT_INIT = 16'he4aa;
    SB_DFF i251_252 (.Q(\mem_LUT.mem_2_7 ), .C(SLM_CLK_c), .D(n6053));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i248_249 (.Q(\mem_LUT.mem_2_6 ), .C(SLM_CLK_c), .D(n6052));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i245_246 (.Q(\mem_LUT.mem_2_5 ), .C(SLM_CLK_c), .D(n6051));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i242_243 (.Q(\mem_LUT.mem_2_4 ), .C(SLM_CLK_c), .D(n6050));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i239_240 (.Q(\mem_LUT.mem_2_3 ), .C(SLM_CLK_c), .D(n6049));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i236_237 (.Q(\mem_LUT.mem_2_2 ), .C(SLM_CLK_c), .D(n6048));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i233_234 (.Q(\mem_LUT.mem_2_1 ), .C(SLM_CLK_c), .D(n6047));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i230_231 (.Q(\mem_LUT.mem_2_0 ), .C(SLM_CLK_c), .D(n6046));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i155_156 (.Q(\mem_LUT.mem_1_7 ), .C(SLM_CLK_c), .D(n6040));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i152_153 (.Q(\mem_LUT.mem_1_6 ), .C(SLM_CLK_c), .D(n6039));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i149_150 (.Q(\mem_LUT.mem_1_5 ), .C(SLM_CLK_c), .D(n6038));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i146_147 (.Q(\mem_LUT.mem_1_4 ), .C(SLM_CLK_c), .D(n6037));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i143_144 (.Q(\mem_LUT.mem_1_3 ), .C(SLM_CLK_c), .D(n6036));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i140_141 (.Q(\mem_LUT.mem_1_2 ), .C(SLM_CLK_c), .D(n6035));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i137_138 (.Q(\mem_LUT.mem_1_1 ), .C(SLM_CLK_c), .D(n6034));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 n12557_bdd_4_lut (.I0(n12557), .I1(\mem_LUT.mem_1_4 ), .I2(\mem_LUT.mem_0_4 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1084 [4]));
    defparam n12557_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i134_135 (.Q(\mem_LUT.mem_1_0 ), .C(SLM_CLK_c), .D(n6033));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i59_60 (.Q(\mem_LUT.mem_0_7 ), .C(SLM_CLK_c), .D(n6032));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i56_57 (.Q(\mem_LUT.mem_0_6 ), .C(SLM_CLK_c), .D(n6031));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i53_54 (.Q(\mem_LUT.mem_0_5 ), .C(SLM_CLK_c), .D(n6030));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i50_51 (.Q(\mem_LUT.mem_0_4 ), .C(SLM_CLK_c), .D(n6029));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i47_48 (.Q(\mem_LUT.mem_0_3 ), .C(SLM_CLK_c), .D(n6028));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i44_45 (.Q(\mem_LUT.mem_0_2 ), .C(SLM_CLK_c), .D(n6027));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i41_42 (.Q(\mem_LUT.mem_0_1 ), .C(SLM_CLK_c), .D(n6026));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i38_39 (.Q(\mem_LUT.mem_0_0 ), .C(SLM_CLK_c), .D(n6025));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 i1394_3_lut (.I0(wr_addr_r[2]), .I1(wr_addr_r[1]), .I2(wr_addr_r[0]), 
            .I3(GND_net), .O(\wr_addr_p1_w[2] ));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam i1394_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1_4_lut (.I0(n1), .I1(\wr_addr_p1_w[2] ), .I2(n2), .I3(rd_addr_r[2]), 
            .O(n10226));
    defparam i1_4_lut.LUT_INIT = 16'h0208;
    SB_LUT4 wr_addr_r_1__I_0_i1_2_lut (.I0(wr_addr_r[0]), .I1(rd_addr_r[0]), 
            .I2(GND_net), .I3(GND_net), .O(n1));   // src/fifo_quad_word_mod.v(115[26:58])
    defparam wr_addr_r_1__I_0_i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE wr_addr_r__i2 (.Q(wr_addr_r[2]), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n5989));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF \mem_LUT.data_buff_r__i4  (.Q(\fifo_temp_output[4] ), .C(SLM_CLK_c), 
           .D(n5311));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i5  (.Q(\fifo_temp_output[5] ), .C(SLM_CLK_c), 
           .D(n5314));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10672 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_3 ), 
            .I2(\mem_LUT.mem_3_3 ), .I3(rd_addr_r[1]), .O(n12491));
    defparam rd_addr_r_0__bdd_4_lut_10672.LUT_INIT = 16'he4aa;
    SB_LUT4 n12491_bdd_4_lut (.I0(n12491), .I1(\mem_LUT.mem_1_3 ), .I2(\mem_LUT.mem_0_3 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1084 [3]));
    defparam n12491_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4685_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_3_7 ), .O(n6068));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4685_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE wr_addr_r__i1 (.Q(wr_addr_r[1]), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n5868));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF \mem_LUT.data_buff_r__i2  (.Q(\fifo_temp_output[2] ), .C(SLM_CLK_c), 
           .D(n4882));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10617 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_2 ), 
            .I2(\mem_LUT.mem_3_2 ), .I3(rd_addr_r[1]), .O(n12485));
    defparam rd_addr_r_0__bdd_4_lut_10617.LUT_INIT = 16'he4aa;
    SB_LUT4 n12485_bdd_4_lut (.I0(n12485), .I1(\mem_LUT.mem_1_2 ), .I2(\mem_LUT.mem_0_2 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1084 [2]));
    defparam n12485_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF \mem_LUT.data_buff_r__i3  (.Q(\fifo_temp_output[3] ), .C(SLM_CLK_c), 
           .D(n4887));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10612 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_1 ), 
            .I2(\mem_LUT.mem_3_1 ), .I3(rd_addr_r[1]), .O(n12473));
    defparam rd_addr_r_0__bdd_4_lut_10612.LUT_INIT = 16'he4aa;
    SB_LUT4 n12473_bdd_4_lut (.I0(n12473), .I1(\mem_LUT.mem_1_1 ), .I2(\mem_LUT.mem_0_1 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1084 [1]));
    defparam n12473_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF \mem_LUT.data_buff_r__i6  (.Q(\fifo_temp_output[6] ), .C(SLM_CLK_c), 
           .D(n5536));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i7  (.Q(\fifo_temp_output[7] ), .C(SLM_CLK_c), 
           .D(n5539));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 i4684_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_3_6 ), .O(n6067));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4684_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF empty_r_85 (.Q(is_fifo_empty_flag), .C(SLM_CLK_c), .D(n10786));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10602 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_0 ), 
            .I2(\mem_LUT.mem_3_0 ), .I3(rd_addr_r[1]), .O(n12437));
    defparam rd_addr_r_0__bdd_4_lut_10602.LUT_INIT = 16'he4aa;
    SB_LUT4 n12437_bdd_4_lut (.I0(n12437), .I1(\mem_LUT.mem_1_0 ), .I2(\mem_LUT.mem_0_0 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1084 [0]));
    defparam n12437_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4683_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_3_5 ), .O(n6066));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4683_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4682_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_3_4 ), .O(n6065));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4682_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF rd_addr_r__i1 (.Q(rd_addr_r[1]), .C(SLM_CLK_c), .D(n4919));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 i4681_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_3_3 ), .O(n6064));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4681_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4680_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_3_2 ), .O(n6063));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4680_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF rd_addr_r__i2 (.Q(rd_addr_r[2]), .C(SLM_CLK_c), .D(n4922));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 i4679_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_3_1 ), .O(n6062));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4679_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4678_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_3_0 ), .O(n6061));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4678_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4670_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_2_7 ), .O(n6053));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4670_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4669_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_2_6 ), .O(n6052));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4669_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4668_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_2_5 ), .O(n6051));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4668_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4667_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_2_4 ), .O(n6050));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4667_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4666_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_2_3 ), .O(n6049));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4666_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4665_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_2_2 ), .O(n6048));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4665_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_en_i_I_0_2_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(GND_net), .I3(GND_net), .O(wr_fifo_en_w));   // src/fifo_quad_word_mod.v(103[21:60])
    defparam wr_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4664_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_2_1 ), .O(n6047));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4664_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4663_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_2_0 ), .O(n6046));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4663_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF rd_fifo_en_prev_r_86 (.Q(rd_fifo_en_prev_r), .C(SLM_CLK_c), .D(n4878));   // src/fifo_quad_word_mod.v(353[29] 363[32])
    SB_LUT4 rd_en_i_I_0_2_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(GND_net), .I3(GND_net), .O(rd_fifo_en_w));   // src/fifo_quad_word_mod.v(62[29:51])
    defparam rd_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4657_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_1_7 ), .O(n6040));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4657_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4656_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_1_6 ), .O(n6039));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4656_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4655_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_1_5 ), .O(n6038));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4655_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4654_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_1_4 ), .O(n6037));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4654_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4653_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_1_3 ), .O(n6036));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4653_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4652_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_1_2 ), .O(n6035));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4652_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4651_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_1_1 ), .O(n6034));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4651_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4650_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_1_0 ), .O(n6033));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4650_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4649_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_0_7 ), .O(n6032));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4649_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4648_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_0_6 ), .O(n6031));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4648_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4647_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_0_5 ), .O(n6030));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4647_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4646_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_0_4 ), .O(n6029));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4646_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4645_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_0_3 ), .O(n6028));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4645_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4644_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_0_2 ), .O(n6027));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4644_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4643_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_0_1 ), .O(n6026));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4643_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4642_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_0_0 ), .O(n6025));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4642_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1603_2_lut_4_lut (.I0(rd_addr_r[0]), .I1(fifo_read_cmd), .I2(is_fifo_empty_flag), 
            .I3(reset_all_w), .O(n12[0]));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1603_2_lut_4_lut.LUT_INIT = 16'h55a6;
    SB_LUT4 EnabledDecoder_2_i3_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(GND_net), .O(n3));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i3_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i4_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(GND_net), .O(n4));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i4_2_lut_3_lut.LUT_INIT = 16'h0202;
    
endmodule
//
// Verilog Description of module spi
//

module spi (\tx_data_byte[3] , n2086, GND_net, \tx_data_byte[4] , SEN_c_1, 
            SLM_CLK_c, \tx_data_byte[5] , SOUT_c, n4312, \rx_shift_reg[0] , 
            \tx_data_byte[6] , n4319, SDAT_c_15, \tx_data_byte[7] , 
            tx_addr_byte, VCC_net, n10428, \tx_shift_reg[0] , n6060, 
            rx_buf_byte, n6059, n6058, n6057, n6056, n6055, n6054, 
            spi_rx_byte_ready, SCK_c_0, spi_start_transfer_r, n4897, 
            n4888, \rx_shift_reg[1] , n4883, \rx_shift_reg[2] , n4877, 
            \rx_shift_reg[3] , n4869, \rx_shift_reg[4] , n4838, \rx_shift_reg[5] , 
            multi_byte_spi_trans_flag_r, n4836, \rx_shift_reg[6] , n4834, 
            \rx_shift_reg[7] , \tx_data_byte[2] , \tx_data_byte[1] , n3495) /* synthesis syn_module_defined=1 */ ;
    input \tx_data_byte[3] ;
    output n2086;
    input GND_net;
    input \tx_data_byte[4] ;
    output SEN_c_1;
    input SLM_CLK_c;
    input \tx_data_byte[5] ;
    input SOUT_c;
    output n4312;
    output \rx_shift_reg[0] ;
    input \tx_data_byte[6] ;
    output n4319;
    output SDAT_c_15;
    input \tx_data_byte[7] ;
    input [7:0]tx_addr_byte;
    input VCC_net;
    input n10428;
    output \tx_shift_reg[0] ;
    input n6060;
    output [7:0]rx_buf_byte;
    input n6059;
    input n6058;
    input n6057;
    input n6056;
    input n6055;
    input n6054;
    output spi_rx_byte_ready;
    output SCK_c_0;
    input spi_start_transfer_r;
    input n4897;
    input n4888;
    output \rx_shift_reg[1] ;
    input n4883;
    output \rx_shift_reg[2] ;
    input n4877;
    output \rx_shift_reg[3] ;
    input n4869;
    output \rx_shift_reg[4] ;
    input n4838;
    output \rx_shift_reg[5] ;
    input multi_byte_spi_trans_flag_r;
    input n4836;
    output \rx_shift_reg[6] ;
    input n4834;
    output \rx_shift_reg[7] ;
    input \tx_data_byte[2] ;
    input \tx_data_byte[1] ;
    output n3495;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [15:0]tx_shift_reg;   // src/spi.v(70[12:24])
    wire [15:0]n2087;
    
    wire n7109;
    wire [3:0]state;   // src/spi.v(71[11:16])
    
    wire n12080;
    wire [9:0]counter;   // src/spi.v(69[11:18])
    
    wire n12081;
    wire [2:0]n970;
    wire [3:0]state_3__N_938;
    
    wire n10827, n24, n12108;
    wire [9:0]n45;
    
    wire n4380, n4694, n10203, n10204, n10202, n10201, n10200, 
        n10199, n10198, n10197, n10196;
    wire [7:0]n315;
    wire [7:0]multi_byte_counter;   // src/spi.v(68[11:29])
    wire [7:0]n2142;
    
    wire n10171, n10170, n10169, n10168, n10167, n10166, n10165, 
        n4, n37, n2, n4_adj_2, n51_adj_3, n12072, n3748, n12073, 
        n14, n19, n12052, n12057, n34, n37_adj_4, n10851, n4236, 
        n19_adj_5, n10778, n7, n4358, n10828, n10792, n10826, 
        n4_adj_6, n4629, n4541, n4672, n10, n14_adj_7, n34_adj_8, 
        n10_adj_9, n14_adj_10, n12101, n7_adj_11, n3, n3_adj_12, 
        n21, n10941, n22, n3_adj_13, n4519, n12112, n7_adj_14, 
        n12104;
    
    SB_LUT4 mux_981_i4_3_lut (.I0(\tx_data_byte[3] ), .I1(tx_shift_reg[2]), 
            .I2(n2086), .I3(GND_net), .O(n2087[3]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i5_3_lut (.I0(\tx_data_byte[4] ), .I1(tx_shift_reg[3]), 
            .I2(n2086), .I3(GND_net), .O(n2087[4]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10320_4_lut (.I0(n7109), .I1(state[1]), .I2(state[0]), .I3(state[2]), 
            .O(n12080));   // src/spi.v(88[9] 219[16])
    defparam i10320_4_lut.LUT_INIT = 16'hc08c;
    SB_LUT4 i1_4_lut (.I0(counter[4]), .I1(n12080), .I2(n12081), .I3(state[3]), 
            .O(n970[0]));   // src/spi.v(76[8] 221[4])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_DFF byte_recv_92_i2 (.Q(SEN_c_1), .C(SLM_CLK_c), .D(n970[1]));   // src/spi.v(88[9] 219[16])
    SB_LUT4 mux_981_i6_3_lut (.I0(\tx_data_byte[5] ), .I1(tx_shift_reg[4]), 
            .I2(n2086), .I3(GND_net), .O(n2087[5]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE rx_shift_reg_i0 (.Q(\rx_shift_reg[0] ), .C(SLM_CLK_c), .E(n4312), 
            .D(SOUT_c));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i0 (.Q(state[0]), .C(SLM_CLK_c), .E(n10827), .D(state_3__N_938[0]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i1_2_lut_3_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(GND_net), .O(n24));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i10319_2_lut_3_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(GND_net), .O(n12108));
    defparam i10319_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFFESR counter_1189__i0 (.Q(counter[0]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[0]), .R(n4694));   // src/spi.v(183[28:41])
    SB_LUT4 mux_981_i7_3_lut (.I0(\tx_data_byte[6] ), .I1(tx_shift_reg[5]), 
            .I2(n2086), .I3(GND_net), .O(n2087[6]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE tx_shift_reg_i0_i15 (.Q(SDAT_c_15), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[15]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_981_i8_3_lut (.I0(\tx_data_byte[7] ), .I1(tx_shift_reg[6]), 
            .I2(n2086), .I3(GND_net), .O(n2087[7]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i9_3_lut (.I0(tx_addr_byte[0]), .I1(tx_shift_reg[7]), 
            .I2(n2086), .I3(GND_net), .O(n2087[8]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i10_3_lut (.I0(tx_addr_byte[1]), .I1(tx_shift_reg[8]), 
            .I2(n2086), .I3(GND_net), .O(n2087[9]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i11_3_lut (.I0(tx_addr_byte[2]), .I1(tx_shift_reg[9]), 
            .I2(n2086), .I3(GND_net), .O(n2087[10]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i12_3_lut (.I0(tx_addr_byte[3]), .I1(tx_shift_reg[10]), 
            .I2(n2086), .I3(GND_net), .O(n2087[11]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i13_3_lut (.I0(tx_addr_byte[4]), .I1(tx_shift_reg[11]), 
            .I2(n2086), .I3(GND_net), .O(n2087[12]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i14_3_lut (.I0(tx_addr_byte[5]), .I1(tx_shift_reg[12]), 
            .I2(n2086), .I3(GND_net), .O(n2087[13]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i15_3_lut (.I0(tx_addr_byte[6]), .I1(tx_shift_reg[13]), 
            .I2(n2086), .I3(GND_net), .O(n2087[14]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY counter_1189_add_4_10 (.CI(n10203), .I0(VCC_net), .I1(counter[8]), 
            .CO(n10204));
    SB_LUT4 counter_1189_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[7]), 
            .I3(n10202), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFE tx_shift_reg_i0_i0 (.Q(\tx_shift_reg[0] ), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n10428));   // src/spi.v(76[8] 221[4])
    SB_CARRY counter_1189_add_4_9 (.CI(n10202), .I0(VCC_net), .I1(counter[7]), 
            .CO(n10203));
    SB_DFF Rx_Recv_Byte_i1 (.Q(rx_buf_byte[1]), .C(SLM_CLK_c), .D(n6060));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i2 (.Q(rx_buf_byte[2]), .C(SLM_CLK_c), .D(n6059));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i3 (.Q(rx_buf_byte[3]), .C(SLM_CLK_c), .D(n6058));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i4 (.Q(rx_buf_byte[4]), .C(SLM_CLK_c), .D(n6057));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i5 (.Q(rx_buf_byte[5]), .C(SLM_CLK_c), .D(n6056));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i6 (.Q(rx_buf_byte[6]), .C(SLM_CLK_c), .D(n6055));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i7 (.Q(rx_buf_byte[7]), .C(SLM_CLK_c), .D(n6054));   // src/spi.v(76[8] 221[4])
    SB_LUT4 counter_1189_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[6]), 
            .I3(n10201), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_8 (.CI(n10201), .I0(VCC_net), .I1(counter[6]), 
            .CO(n10202));
    SB_LUT4 counter_1189_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[5]), 
            .I3(n10200), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_7 (.CI(n10200), .I0(VCC_net), .I1(counter[5]), 
            .CO(n10201));
    SB_LUT4 counter_1189_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[4]), 
            .I3(n10199), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_6 (.CI(n10199), .I0(VCC_net), .I1(counter[4]), 
            .CO(n10200));
    SB_LUT4 counter_1189_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[3]), 
            .I3(n10198), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_5 (.CI(n10198), .I0(VCC_net), .I1(counter[3]), 
            .CO(n10199));
    SB_LUT4 counter_1189_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[2]), 
            .I3(n10197), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_4 (.CI(n10197), .I0(VCC_net), .I1(counter[2]), 
            .CO(n10198));
    SB_LUT4 counter_1189_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[1]), 
            .I3(n10196), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_3 (.CI(n10196), .I0(VCC_net), .I1(counter[1]), 
            .CO(n10197));
    SB_LUT4 counter_1189_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n10196));
    SB_LUT4 add_995_9_lut (.I0(GND_net), .I1(multi_byte_counter[7]), .I2(n2142[5]), 
            .I3(n10171), .O(n315[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_995_8_lut (.I0(GND_net), .I1(multi_byte_counter[6]), .I2(n2142[5]), 
            .I3(n10170), .O(n315[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_8 (.CI(n10170), .I0(multi_byte_counter[6]), .I1(n2142[5]), 
            .CO(n10171));
    SB_LUT4 add_995_7_lut (.I0(GND_net), .I1(multi_byte_counter[5]), .I2(n2142[5]), 
            .I3(n10169), .O(n315[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_7 (.CI(n10169), .I0(multi_byte_counter[5]), .I1(n2142[5]), 
            .CO(n10170));
    SB_LUT4 add_995_6_lut (.I0(GND_net), .I1(multi_byte_counter[4]), .I2(n2142[5]), 
            .I3(n10168), .O(n315[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_6 (.CI(n10168), .I0(multi_byte_counter[4]), .I1(n2142[5]), 
            .CO(n10169));
    SB_LUT4 add_995_5_lut (.I0(GND_net), .I1(multi_byte_counter[3]), .I2(n2142[5]), 
            .I3(n10167), .O(n315[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_5 (.CI(n10167), .I0(multi_byte_counter[3]), .I1(n2142[5]), 
            .CO(n10168));
    SB_LUT4 add_995_4_lut (.I0(GND_net), .I1(multi_byte_counter[2]), .I2(n2142[5]), 
            .I3(n10166), .O(n315[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_4 (.CI(n10166), .I0(multi_byte_counter[2]), .I1(n2142[5]), 
            .CO(n10167));
    SB_LUT4 add_995_3_lut (.I0(GND_net), .I1(multi_byte_counter[1]), .I2(n2142[5]), 
            .I3(n10165), .O(n315[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_3 (.CI(n10165), .I0(multi_byte_counter[1]), .I1(n2142[5]), 
            .CO(n10166));
    SB_LUT4 add_995_2_lut (.I0(GND_net), .I1(multi_byte_counter[0]), .I2(n2142[5]), 
            .I3(GND_net), .O(n315[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_2 (.CI(GND_net), .I0(multi_byte_counter[0]), .I1(n2142[5]), 
            .CO(n10165));
    SB_DFFE tx_shift_reg_i0_i14 (.Q(tx_shift_reg[14]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[14]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i13 (.Q(tx_shift_reg[13]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[13]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i12 (.Q(tx_shift_reg[12]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[12]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i11 (.Q(tx_shift_reg[11]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[11]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i10 (.Q(tx_shift_reg[10]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[10]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i9 (.Q(tx_shift_reg[9]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[9]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i8 (.Q(tx_shift_reg[8]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[8]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i7 (.Q(tx_shift_reg[7]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[7]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i6 (.Q(tx_shift_reg[6]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[6]));   // src/spi.v(76[8] 221[4])
    SB_DFF byte_recv_92_i3 (.Q(spi_rx_byte_ready), .C(SLM_CLK_c), .D(n970[2]));   // src/spi.v(88[9] 219[16])
    SB_DFFE tx_shift_reg_i0_i5 (.Q(tx_shift_reg[5]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[5]));   // src/spi.v(76[8] 221[4])
    SB_DFF byte_recv_92_i1 (.Q(SCK_c_0), .C(SLM_CLK_c), .D(n970[0]));   // src/spi.v(88[9] 219[16])
    SB_DFFE tx_shift_reg_i0_i4 (.Q(tx_shift_reg[4]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[4]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i3 (.Q(tx_shift_reg[3]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[3]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i1_2_lut (.I0(state[3]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n4));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_3 (.I0(n37), .I1(state[0]), .I2(n2), .I3(n4_adj_2), 
            .O(n2086));
    defparam i1_4_lut_adj_3.LUT_INIT = 16'ha2a0;
    SB_LUT4 i1_2_lut_adj_4 (.I0(counter[4]), .I1(n51_adj_3), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // src/spi.v(183[28:41])
    defparam i1_2_lut_adj_4.LUT_INIT = 16'h4444;
    SB_LUT4 i10314_4_lut (.I0(spi_start_transfer_r), .I1(state[0]), .I2(n37), 
            .I3(state[3]), .O(n12072));   // src/spi.v(71[11:16])
    defparam i10314_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1_4_lut_adj_5 (.I0(n3748), .I1(n12072), .I2(n12073), .I3(state[1]), 
            .O(n4319));
    defparam i1_4_lut_adj_5.LUT_INIT = 16'h5044;
    SB_LUT4 mux_981_i16_3_lut (.I0(tx_addr_byte[7]), .I1(tx_shift_reg[14]), 
            .I2(n2086), .I3(GND_net), .O(n2087[15]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(state[3]), .I1(state[2]), .I2(state[0]), .I3(GND_net), 
            .O(n14));   // src/spi.v(88[9] 219[16])
    defparam i1_3_lut.LUT_INIT = 16'hcdcd;
    SB_LUT4 i10301_3_lut (.I0(state[0]), .I1(state[2]), .I2(n19), .I3(GND_net), 
            .O(n12052));
    defparam i10301_3_lut.LUT_INIT = 16'h4d4d;
    SB_LUT4 i10298_3_lut (.I0(state[3]), .I1(state[2]), .I2(state[0]), 
            .I3(GND_net), .O(n12057));
    defparam i10298_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF Rx_Recv_Byte_i0 (.Q(rx_buf_byte[0]), .C(SLM_CLK_c), .D(n4897));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i65_3_lut (.I0(n14), .I1(n12052), .I2(state[1]), .I3(GND_net), 
            .O(n34));
    defparam i65_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i66_4_lut (.I0(n12057), .I1(n2142[5]), .I2(state[1]), .I3(state[3]), 
            .O(n37_adj_4));
    defparam i66_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_4_lut_adj_6 (.I0(state[3]), .I1(n37_adj_4), .I2(n34), .I3(n10851), 
            .O(n4694));
    defparam i1_4_lut_adj_6.LUT_INIT = 16'h50dc;
    SB_LUT4 i10430_4_lut (.I0(state[3]), .I1(state[1]), .I2(n4236), .I3(n14), 
            .O(n4380));   // src/spi.v(88[9] 219[16])
    defparam i10430_4_lut.LUT_INIT = 16'h4c5f;
    SB_DFF rx_shift_reg_i1 (.Q(\rx_shift_reg[1] ), .C(SLM_CLK_c), .D(n4888));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i2 (.Q(tx_shift_reg[2]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[2]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i1 (.Q(tx_shift_reg[1]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[1]));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i2 (.Q(\rx_shift_reg[2] ), .C(SLM_CLK_c), .D(n4883));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i3 (.Q(state[3]), .C(SLM_CLK_c), .E(n19_adj_5), .D(state_3__N_938[3]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i2_3_lut (.I0(state[3]), .I1(n19), .I2(state[1]), .I3(GND_net), 
            .O(n10778));
    defparam i2_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i4_4_lut (.I0(n7), .I1(state[3]), .I2(spi_start_transfer_r), 
            .I3(state[0]), .O(n4358));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(state[1]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n7));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFFE state_i2 (.Q(state[2]), .C(SLM_CLK_c), .E(n10828), .D(state_3__N_938[2]));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i1 (.Q(state[1]), .C(SLM_CLK_c), .E(n10792), .D(state_3__N_938[1]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i1_4_lut_adj_7 (.I0(n4358), .I1(n10778), .I2(state[0]), .I3(state[2]), 
            .O(n10826));
    defparam i1_4_lut_adj_7.LUT_INIT = 16'h8aaa;
    SB_DFF rx_shift_reg_i3 (.Q(\rx_shift_reg[3] ), .C(SLM_CLK_c), .D(n4877));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i1_2_lut_adj_8 (.I0(n19), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_6));
    defparam i1_2_lut_adj_8.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_4_lut_adj_9 (.I0(state[3]), .I1(n10826), .I2(n7), .I3(n4_adj_6), 
            .O(n10827));
    defparam i1_4_lut_adj_9.LUT_INIT = 16'h4c44;
    SB_LUT4 i3_4_lut (.I0(counter[0]), .I1(counter[3]), .I2(counter[2]), 
            .I3(counter[1]), .O(n51_adj_3));   // src/spi.v(183[28:41])
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i9015_2_lut (.I0(state[0]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n10851));
    defparam i9015_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_10 (.I0(state[2]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n3748));   // src/spi.v(88[9] 219[16])
    defparam i1_2_lut_adj_10.LUT_INIT = 16'h2222;
    SB_LUT4 i10440_3_lut (.I0(counter[4]), .I1(n4629), .I2(n51_adj_3), 
            .I3(GND_net), .O(n4312));   // src/spi.v(88[9] 219[16])
    defparam i10440_3_lut.LUT_INIT = 16'h2020;
    SB_DFFESR counter_1189__i1 (.Q(counter[1]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[1]), .R(n4694));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1189__i2 (.Q(counter[2]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[2]), .R(n4694));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1189__i3 (.Q(counter[3]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[3]), .R(n4694));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1189__i4 (.Q(counter[4]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[4]), .R(n4694));   // src/spi.v(183[28:41])
    SB_DFF rx_shift_reg_i4 (.Q(\rx_shift_reg[4] ), .C(SLM_CLK_c), .D(n4869));   // src/spi.v(76[8] 221[4])
    SB_DFFESR counter_1189__i5 (.Q(counter[5]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[5]), .R(n4694));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1189__i9 (.Q(counter[9]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[9]), .R(n4694));   // src/spi.v(183[28:41])
    SB_DFFESS counter_1189__i8 (.Q(counter[8]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[8]), .S(n4694));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1189__i7 (.Q(counter[7]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[7]), .R(n4694));   // src/spi.v(183[28:41])
    SB_DFFESR multi_byte_counter_i1 (.Q(multi_byte_counter[1]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[1]), .R(n4672));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i2 (.Q(multi_byte_counter[2]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[2]), .R(n4672));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i3 (.Q(multi_byte_counter[3]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[3]), .R(n4672));   // src/spi.v(76[8] 221[4])
    SB_DFFESR counter_1189__i6 (.Q(counter[6]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[6]), .R(n4694));   // src/spi.v(183[28:41])
    SB_DFFESR multi_byte_counter_i4 (.Q(multi_byte_counter[4]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[4]), .R(n4672));   // src/spi.v(76[8] 221[4])
    SB_DFFESS multi_byte_counter_i5 (.Q(multi_byte_counter[5]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[5]), .S(n4672));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i2_2_lut_adj_11 (.I0(multi_byte_counter[2]), .I1(multi_byte_counter[4]), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // src/spi.v(208[21:52])
    defparam i2_2_lut_adj_11.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(multi_byte_counter[3]), .I1(multi_byte_counter[1]), 
            .I2(multi_byte_counter[5]), .I3(multi_byte_counter[7]), .O(n14_adj_7));   // src/spi.v(208[21:52])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(multi_byte_counter[0]), .I1(n14_adj_7), .I2(n10), 
            .I3(multi_byte_counter[6]), .O(n2142[5]));   // src/spi.v(208[21:52])
    defparam i7_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i2_3_lut_adj_12 (.I0(counter[2]), .I1(counter[1]), .I2(counter[3]), 
            .I3(GND_net), .O(n34_adj_8));   // src/spi.v(183[28:41])
    defparam i2_3_lut_adj_12.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_2_lut_adj_13 (.I0(counter[6]), .I1(counter[7]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_9));   // src/spi.v(141[21:41])
    defparam i2_2_lut_adj_13.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_14 (.I0(counter[4]), .I1(counter[5]), .I2(counter[9]), 
            .I3(n34_adj_8), .O(n14_adj_10));   // src/spi.v(141[21:41])
    defparam i6_4_lut_adj_14.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_15 (.I0(counter[0]), .I1(n14_adj_10), .I2(n10_adj_9), 
            .I3(counter[8]), .O(n19));   // src/spi.v(141[21:41])
    defparam i7_4_lut_adj_15.LUT_INIT = 16'hfffd;
    SB_LUT4 i10345_3_lut (.I0(n2142[5]), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n12101));   // src/spi.v(88[9] 219[16])
    defparam i10345_3_lut.LUT_INIT = 16'hc4c4;
    SB_LUT4 mux_344_Mux_1_i7_4_lut (.I0(state[0]), .I1(state[2]), .I2(n19), 
            .I3(state[1]), .O(n7_adj_11));   // src/spi.v(88[9] 219[16])
    defparam mux_344_Mux_1_i7_4_lut.LUT_INIT = 16'h02dd;
    SB_LUT4 mux_344_Mux_1_i15_4_lut (.I0(n7_adj_11), .I1(n12101), .I2(state[3]), 
            .I3(state[2]), .O(n970[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_344_Mux_1_i15_4_lut.LUT_INIT = 16'hfaca;
    SB_DFFESR multi_byte_counter_i0 (.Q(multi_byte_counter[0]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[0]), .R(n4672));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i6 (.Q(multi_byte_counter[6]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[6]), .R(n4672));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i5 (.Q(\rx_shift_reg[5] ), .C(SLM_CLK_c), .D(n4838));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_56_Mux_1_i3_3_lut_3_lut (.I0(multi_byte_spi_trans_flag_r), 
            .I1(state[0]), .I2(state[1]), .I3(GND_net), .O(n3));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_1_i3_3_lut_3_lut.LUT_INIT = 16'h3e3e;
    SB_LUT4 mux_56_Mux_0_i3_4_lut_4_lut (.I0(multi_byte_spi_trans_flag_r), 
            .I1(state[0]), .I2(state[1]), .I3(n19), .O(n3_adj_12));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_0_i3_4_lut_4_lut.LUT_INIT = 16'hc131;
    SB_DFFESS multi_byte_counter_i7 (.Q(multi_byte_counter[7]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[7]), .S(n4672));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i6 (.Q(\rx_shift_reg[6] ), .C(SLM_CLK_c), .D(n4836));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i43_4_lut_4_lut (.I0(state[3]), .I1(state[2]), .I2(state[1]), 
            .I3(state[0]), .O(n21));
    defparam i43_4_lut_4_lut.LUT_INIT = 16'hf01a;
    SB_LUT4 i3273_3_lut_4_lut (.I0(state[3]), .I1(state[2]), .I2(state[0]), 
            .I3(n3_adj_12), .O(state_3__N_938[0]));
    defparam i3273_3_lut_4_lut.LUT_INIT = 16'h1f0e;
    SB_DFF rx_shift_reg_i7 (.Q(\rx_shift_reg[7] ), .C(SLM_CLK_c), .D(n4834));   // src/spi.v(76[8] 221[4])
    SB_LUT4 counter_1189_add_4_11_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[9]), 
            .I3(n10204), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1189_add_4_10_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[8]), 
            .I3(n10203), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_981_i3_3_lut (.I0(\tx_data_byte[2] ), .I1(tx_shift_reg[1]), 
            .I2(n2086), .I3(GND_net), .O(n2087[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i2_3_lut (.I0(\tx_data_byte[1] ), .I1(\tx_shift_reg[0] ), 
            .I2(n2086), .I3(GND_net), .O(n2087[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[2]), .I1(n10778), .I2(n4358), .I3(state[0]), 
            .O(n10828));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hc0e0;
    SB_LUT4 i9104_3_lut_4_lut (.I0(state[0]), .I1(state[2]), .I2(spi_start_transfer_r), 
            .I3(state[1]), .O(n10941));
    defparam i9104_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_56_Mux_3_i15_4_lut (.I0(n12108), .I1(state[1]), .I2(state[3]), 
            .I3(n2142[5]), .O(state_3__N_938[3]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_3_i15_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i10427_4_lut (.I0(n22), .I1(n10941), .I2(n24), .I3(state[3]), 
            .O(n19_adj_5));
    defparam i10427_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i1_2_lut_adj_16 (.I0(n19), .I1(n21), .I2(GND_net), .I3(GND_net), 
            .O(n22));
    defparam i1_2_lut_adj_16.LUT_INIT = 16'h8888;
    SB_LUT4 i10306_2_lut_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(n7109), .O(n12081));   // src/spi.v(88[9] 219[16])
    defparam i10306_2_lut_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 mux_56_Mux_2_i15_4_lut (.I0(n3_adj_13), .I1(state[2]), .I2(state[3]), 
            .I3(state[0]), .O(state_3__N_938[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_2_i15_4_lut.LUT_INIT = 16'hc2ce;
    SB_LUT4 mux_56_Mux_2_i3_3_lut (.I0(multi_byte_spi_trans_flag_r), .I1(state[0]), 
            .I2(state[1]), .I3(GND_net), .O(n3_adj_13));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_2_i3_3_lut.LUT_INIT = 16'hc2c2;
    SB_LUT4 i1_2_lut_adj_17 (.I0(state[2]), .I1(n10778), .I2(GND_net), 
            .I3(GND_net), .O(n4519));
    defparam i1_2_lut_adj_17.LUT_INIT = 16'heeee;
    SB_LUT4 mux_56_Mux_1_i7_4_lut (.I0(n3), .I1(n12112), .I2(state[2]), 
            .I3(state[1]), .O(n7_adj_14));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_1_i7_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i2050_4_lut_4_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(state[3]), .O(n4629));   // src/spi.v(88[9] 219[16])
    defparam i2050_4_lut_4_lut_4_lut.LUT_INIT = 16'hfe75;
    SB_LUT4 i10352_2_lut (.I0(n19), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n12112));   // src/spi.v(88[9] 219[16])
    defparam i10352_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_4_lut (.I0(state[3]), .I1(n4519), .I2(n24), .I3(n4358), 
            .O(n10792));
    defparam i2_4_lut.LUT_INIT = 16'h4c00;
    SB_LUT4 i1_4_lut_adj_18 (.I0(state[1]), .I1(n4), .I2(n12104), .I3(state[0]), 
            .O(n4541));
    defparam i1_4_lut_adj_18.LUT_INIT = 16'ha088;
    SB_LUT4 i10290_3_lut (.I0(state[3]), .I1(state[2]), .I2(n19), .I3(GND_net), 
            .O(n12104));
    defparam i10290_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i3289_2_lut (.I0(n4541), .I1(state[3]), .I2(GND_net), .I3(GND_net), 
            .O(n4672));   // src/spi.v(76[8] 221[4])
    defparam i3289_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_4_lut (.I0(n2142[5]), .I1(state[0]), .I2(state[2]), 
            .I3(state[1]), .O(n4236));   // src/spi.v(88[9] 219[16])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[0]), .I1(state[2]), .I2(state[1]), 
            .I3(state[3]), .O(n2));   // src/spi.v(88[9] 219[16])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h00b0;
    SB_LUT4 i10326_2_lut_3_lut (.I0(counter[4]), .I1(n51_adj_3), .I2(state[3]), 
            .I3(GND_net), .O(n12073));   // src/spi.v(71[11:16])
    defparam i10326_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_3_lut_adj_19 (.I0(state[1]), .I1(state[3]), .I2(state[2]), 
            .I3(GND_net), .O(n4_adj_2));
    defparam i1_2_lut_3_lut_adj_19.LUT_INIT = 16'h0404;
    SB_LUT4 i2123_4_lut_4_lut (.I0(state[0]), .I1(state[2]), .I2(state[1]), 
            .I3(state[3]), .O(n3495));   // src/spi.v(88[9] 219[16])
    defparam i2123_4_lut_4_lut.LUT_INIT = 16'hfdfb;
    SB_LUT4 mux_344_Mux_2_i15_4_lut_4_lut (.I0(state[0]), .I1(state[1]), 
            .I2(state[2]), .I3(state[3]), .O(n970[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_344_Mux_2_i15_4_lut_4_lut.LUT_INIT = 16'h0420;
    SB_LUT4 mux_56_Mux_1_i15_3_lut_4_lut (.I0(state[0]), .I1(state[1]), 
            .I2(state[3]), .I3(n7_adj_14), .O(state_3__N_938[1]));
    defparam mux_56_Mux_1_i15_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i1_2_lut_4_lut_adj_20 (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(counter[3]), .O(n7109));   // src/spi.v(183[28:41])
    defparam i1_2_lut_4_lut_adj_20.LUT_INIT = 16'hfffe;
    
endmodule
//
// Verilog Description of module \uart_tx(CLKS_PER_BIT=20) 
//

module \uart_tx(CLKS_PER_BIT=20)  (UART_TX_c, SLM_CLK_c, r_SM_Main, GND_net, 
            \r_SM_Main_2__N_841[1] , \r_SM_Main_2__N_844[0] , n3794, VCC_net, 
            n13865, n10805, n4890, r_Tx_Data, n4889, tx_uart_active_flag, 
            n5192, n5191, n5190, n5189, n5187, n5171, n5170) /* synthesis syn_module_defined=1 */ ;
    output UART_TX_c;
    input SLM_CLK_c;
    output [2:0]r_SM_Main;
    input GND_net;
    output \r_SM_Main_2__N_841[1] ;
    input \r_SM_Main_2__N_844[0] ;
    output n3794;
    input VCC_net;
    input n13865;
    output n10805;
    input n4890;
    output [7:0]r_Tx_Data;
    input n4889;
    output tx_uart_active_flag;
    input n5192;
    input n5191;
    input n5190;
    input n5189;
    input n5187;
    input n5171;
    input n5170;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n3, n1, n3063;
    wire [9:0]n45;
    wire [9:0]r_Clock_Count;   // src/uart_tx.v(32[16:29])
    
    wire n4797, n7576, n10955, n10961;
    wire [2:0]r_Bit_Index;   // src/uart_tx.v(33[16:27])
    
    wire n6098, n3_adj_1, n10222, n10221, n10220, n10219, n10218, 
        n10217, n10216, n10215, n10214;
    wire [2:0]n312;
    
    wire n4, n8, n7, n3062, o_Tx_Serial_N_873, n11099, n11100, 
        n12803, n11082, n11081;
    
    SB_DFFE o_Tx_Serial_44 (.Q(UART_TX_c), .C(SLM_CLK_c), .E(n1), .D(n3));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(SLM_CLK_c), .D(n3063), 
            .R(r_SM_Main[2]));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Clock_Count_1193__i0 (.Q(r_Clock_Count[0]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[0]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_LUT4 i10402_2_lut_3_lut (.I0(n7576), .I1(r_SM_Main[1]), .I2(n10955), 
            .I3(GND_net), .O(n10961));   // src/uart_tx.v(41[7] 140[14])
    defparam i10402_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i4715_3_lut_4_lut (.I0(n7576), .I1(r_SM_Main[1]), .I2(r_Bit_Index[0]), 
            .I3(n10955), .O(n6098));   // src/uart_tx.v(41[7] 140[14])
    defparam i4715_3_lut_4_lut.LUT_INIT = 16'h04f0;
    SB_LUT4 i10400_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_841[1] ), .O(n10955));
    defparam i10400_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_844[0] ), .O(n3794));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n6098));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(SLM_CLK_c), .D(n13865));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(SLM_CLK_c), .D(n3_adj_1), 
            .R(r_SM_Main[2]));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 r_Clock_Count_1193_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[9]), .I3(n10222), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1193_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n10221), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_10 (.CI(n10221), .I0(GND_net), .I1(r_Clock_Count[8]), 
            .CO(n10222));
    SB_LUT4 r_Clock_Count_1193_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n10220), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_9 (.CI(n10220), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n10221));
    SB_LUT4 r_Clock_Count_1193_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n10219), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_8 (.CI(n10219), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n10220));
    SB_LUT4 r_Clock_Count_1193_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n10218), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_7 (.CI(n10218), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n10219));
    SB_LUT4 r_Clock_Count_1193_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n10217), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_6 (.CI(n10217), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n10218));
    SB_LUT4 r_Clock_Count_1193_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n10216), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_5 (.CI(n10216), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n10217));
    SB_LUT4 r_Clock_Count_1193_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n10215), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_4 (.CI(n10215), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n10216));
    SB_LUT4 r_Clock_Count_1193_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n10214), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_3 (.CI(n10214), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n10215));
    SB_LUT4 r_Clock_Count_1193_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n10214));
    SB_DFFESR r_Clock_Count_1193__i9 (.Q(r_Clock_Count[9]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[9]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i8 (.Q(r_Clock_Count[8]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[8]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i7 (.Q(r_Clock_Count[7]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[7]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i6 (.Q(r_Clock_Count[6]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[6]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i5 (.Q(r_Clock_Count[5]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[5]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i4 (.Q(r_Clock_Count[4]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[4]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i3 (.Q(r_Clock_Count[3]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[3]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i2 (.Q(r_Clock_Count[2]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[2]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i1 (.Q(r_Clock_Count[1]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[1]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_LUT4 i10362_4_lut_4_lut (.I0(\r_SM_Main_2__N_841[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_844[0] ), .O(n10805));
    defparam i10362_4_lut_4_lut.LUT_INIT = 16'h8380;
    SB_LUT4 i2385_2_lut_3_lut (.I0(\r_SM_Main_2__N_841[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_1));
    defparam i2385_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_DFF r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(SLM_CLK_c), .D(n4890));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Active_46 (.Q(tx_uart_active_flag), .C(SLM_CLK_c), .D(n4889));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(SLM_CLK_c), .D(n5192));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(SLM_CLK_c), .D(n5191));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(SLM_CLK_c), .D(n5190));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(SLM_CLK_c), .D(n5189));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(SLM_CLK_c), .D(n5187));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i10392_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_841[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n4797));
    defparam i10392_4_lut.LUT_INIT = 16'h4445;
    SB_DFF r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(SLM_CLK_c), .D(n5171));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(SLM_CLK_c), .D(n5170));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(SLM_CLK_c), .E(n10955), 
            .D(n312[1]), .R(n10961));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(SLM_CLK_c), .E(n10955), 
            .D(n312[2]), .R(n10961));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i1_3_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[1]), 
            .I3(GND_net), .O(n4));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i2_2_lut (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[9]), .I2(GND_net), 
            .I3(GND_net), .O(n8));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[6]), .I2(r_Clock_Count[4]), 
            .I3(n4), .O(n7));
    defparam i1_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i5_4_lut (.I0(r_Clock_Count[5]), .I1(n7), .I2(r_Clock_Count[8]), 
            .I3(n8), .O(\r_SM_Main_2__N_841[1] ));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1694_4_lut (.I0(\r_SM_Main_2__N_844[0] ), .I1(n7576), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_841[1] ), .O(n3062));   // src/uart_tx.v(41[7] 140[14])
    defparam i1694_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1695_3_lut (.I0(n3062), .I1(\r_SM_Main_2__N_841[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n3063));   // src/uart_tx.v(41[7] 140[14])
    defparam i1695_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1372_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n312[2]));
    defparam i1372_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 r_SM_Main_2__I_0_55_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_873), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // src/uart_tx.v(41[7] 140[14])
    defparam r_SM_Main_2__I_0_55_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(n7576));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n11099), 
            .I2(n11100), .I3(r_Bit_Index[2]), .O(n12803));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n12803_bdd_4_lut (.I0(n12803), .I1(n11082), .I2(n11081), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_873));
    defparam n12803_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1365_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n312[1]));   // src/uart_tx.v(96[36:51])
    defparam i1365_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9261_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n11099));
    defparam i9261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9262_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n11100));
    defparam i9262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9244_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n11082));
    defparam i9244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9243_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n11081));
    defparam i9243_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module usb3_if
//

module usb3_if (reset_per_frame, reset_per_frame_latched, SLM_CLK_c, DEBUG_3_c, 
            DEBUG_2_c, FIFO_CLK_c, \dc32_fifo_data_in[0] , DEBUG_5_c, 
            buffer_switch_done, buffer_switch_done_latched, VCC_net, FT_OE_c, 
            n571, GND_net, n575, write_to_dc32_fifo_latched_N_425, n2352, 
            n4911, n4910, n4907, FIFO_D15_c_15, FIFO_D14_c_14, FIFO_D13_c_13, 
            FIFO_D12_c_12, FIFO_D11_c_11, FIFO_D10_c_10, FIFO_D9_c_9, 
            FIFO_D8_c_8, FIFO_D7_c_7, FIFO_D6_c_6, FIFO_D5_c_5, FIFO_D4_c_4, 
            FIFO_D3_c_3, FIFO_D2_c_2, FIFO_D1_c_1, dc32_fifo_almost_full, 
            \dc32_fifo_data_in[15] , \dc32_fifo_data_in[14] , \dc32_fifo_data_in[13] , 
            \dc32_fifo_data_in[12] , \dc32_fifo_data_in[11] , \dc32_fifo_data_in[10] , 
            \dc32_fifo_data_in[9] , \dc32_fifo_data_in[8] , \dc32_fifo_data_in[7] , 
            \dc32_fifo_data_in[6] , \dc32_fifo_data_in[5] , \dc32_fifo_data_in[4] , 
            \dc32_fifo_data_in[3] , \dc32_fifo_data_in[2] , \dc32_fifo_data_in[1] , 
            DEBUG_1_c_c, FT_OE_N_420) /* synthesis syn_module_defined=1 */ ;
    input reset_per_frame;
    output reset_per_frame_latched;
    input SLM_CLK_c;
    input DEBUG_3_c;
    output DEBUG_2_c;
    input FIFO_CLK_c;
    output \dc32_fifo_data_in[0] ;
    output DEBUG_5_c;
    input buffer_switch_done;
    output buffer_switch_done_latched;
    input VCC_net;
    output FT_OE_c;
    output n571;
    input GND_net;
    output n575;
    input write_to_dc32_fifo_latched_N_425;
    output n2352;
    input n4911;
    input n4910;
    input n4907;
    input FIFO_D15_c_15;
    input FIFO_D14_c_14;
    input FIFO_D13_c_13;
    input FIFO_D12_c_12;
    input FIFO_D11_c_11;
    input FIFO_D10_c_10;
    input FIFO_D9_c_9;
    input FIFO_D8_c_8;
    input FIFO_D7_c_7;
    input FIFO_D6_c_6;
    input FIFO_D5_c_5;
    input FIFO_D4_c_4;
    input FIFO_D3_c_3;
    input FIFO_D2_c_2;
    input FIFO_D1_c_1;
    input dc32_fifo_almost_full;
    output \dc32_fifo_data_in[15] ;
    output \dc32_fifo_data_in[14] ;
    output \dc32_fifo_data_in[13] ;
    output \dc32_fifo_data_in[12] ;
    output \dc32_fifo_data_in[11] ;
    output \dc32_fifo_data_in[10] ;
    output \dc32_fifo_data_in[9] ;
    output \dc32_fifo_data_in[8] ;
    output \dc32_fifo_data_in[7] ;
    output \dc32_fifo_data_in[6] ;
    output \dc32_fifo_data_in[5] ;
    output \dc32_fifo_data_in[4] ;
    output \dc32_fifo_data_in[3] ;
    output \dc32_fifo_data_in[2] ;
    output \dc32_fifo_data_in[1] ;
    input DEBUG_1_c_c;
    input FT_OE_N_420;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    
    wire dc32_fifo_empty_latched, FT_RD_N_422;
    wire [31:0]dc32_fifo_data_in_latched;   // src/usb3_if.v(68[12:37])
    
    wire write_to_dc32_fifo_latched, FT_OE_N_419, n3004;
    wire [15:0]n562;
    
    wire n618, n3002;
    wire [3:0]state_timeout_counter;   // src/usb3_if.v(66[11:32])
    
    wire n3942, n3014, n3938, n524, n606, n2415, n2408, n608, 
        n2992, n10282, n613;
    wire [10:0]num_lines_clocked_out_10__N_371;
    wire [10:0]num_lines_clocked_out;   // src/usb3_if.v(65[12:33])
    
    wire n10155, n10156;
    wire [10:0]n1;
    
    wire n10164, n10163, n10162, n10161, n10160, n10159, n10158, 
        n10157, n520, n551, n4, n21, n4224, n2400, n4310, n4688, 
        n18, n2401, n16, n20, n2402, n522, n2983, n4181, n4486, 
        n2399, n2390, n3940, n10783, n2266, n12077, n12030;
    
    SB_DFF reset_per_frame_latched_89 (.Q(reset_per_frame_latched), .C(SLM_CLK_c), 
           .D(reset_per_frame));   // src/usb3_if.v(72[8] 85[4])
    SB_DFF dc32_fifo_empty_latched_90 (.Q(dc32_fifo_empty_latched), .C(SLM_CLK_c), 
           .D(DEBUG_3_c));   // src/usb3_if.v(72[8] 85[4])
    SB_DFFSS FT_RD_92 (.Q(DEBUG_2_c), .C(FIFO_CLK_c), .D(FT_RD_N_422), 
            .S(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFN dc32_fifo_data_in_i1 (.Q(\dc32_fifo_data_in[0] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[0]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN write_to_dc32_fifo_99 (.Q(DEBUG_5_c), .C(FIFO_CLK_c), .D(write_to_dc32_fifo_latched));   // src/usb3_if.v(194[8] 197[4])
    SB_DFF buffer_switch_done_latched_88 (.Q(buffer_switch_done_latched), 
           .C(SLM_CLK_c), .D(buffer_switch_done));   // src/usb3_if.v(72[8] 85[4])
    SB_DFFESS FT_OE_91 (.Q(FT_OE_c), .C(FIFO_CLK_c), .E(VCC_net), .D(FT_OE_N_419), 
            .S(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFSS state_FSM_i1 (.Q(n562[0]), .C(FIFO_CLK_c), .D(n3004), .S(reset_per_frame_latched));   // src/usb3_if.v(98[9] 189[16])
    SB_DFFSR state_FSM_i8 (.Q(n571), .C(FIFO_CLK_c), .D(n618), .R(reset_per_frame_latched));   // src/usb3_if.v(98[9] 189[16])
    SB_DFFSR state_FSM_i7 (.Q(n562[6]), .C(FIFO_CLK_c), .D(n3002), .R(reset_per_frame_latched));   // src/usb3_if.v(98[9] 189[16])
    SB_LUT4 i1_3_lut_4_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[0]), 
            .I2(state_timeout_counter[2]), .I3(state_timeout_counter[3]), 
            .O(n3942));   // src/usb3_if.v(150[42:69])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h01fe;
    SB_DFFSR state_FSM_i6 (.Q(n562[5]), .C(FIFO_CLK_c), .D(n3014), .R(reset_per_frame_latched));   // src/usb3_if.v(98[9] 189[16])
    SB_LUT4 i1_2_lut_3_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[0]), 
            .I2(state_timeout_counter[2]), .I3(GND_net), .O(n3938));   // src/usb3_if.v(150[42:69])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h1e1e;
    SB_LUT4 i1600_3_lut_4_lut (.I0(n562[2]), .I1(n562[0]), .I2(n524), 
            .I3(n606), .O(n2415));   // src/usb3_if.v(98[9] 189[16])
    defparam i1600_3_lut_4_lut.LUT_INIT = 16'h20fd;
    SB_LUT4 i1166_2_lut_3_lut (.I0(n562[2]), .I1(n562[0]), .I2(n524), 
            .I3(GND_net), .O(n2408));   // src/usb3_if.v(98[9] 189[16])
    defparam i1166_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_DFFSR state_FSM_i4 (.Q(n575), .C(FIFO_CLK_c), .D(n608), .R(reset_per_frame_latched));   // src/usb3_if.v(98[9] 189[16])
    SB_DFFSR state_FSM_i3 (.Q(n562[2]), .C(FIFO_CLK_c), .D(n2992), .R(reset_per_frame_latched));   // src/usb3_if.v(98[9] 189[16])
    SB_DFFSR state_FSM_i2 (.Q(n562[1]), .C(FIFO_CLK_c), .D(n10282), .R(reset_per_frame_latched));   // src/usb3_if.v(98[9] 189[16])
    SB_LUT4 i1116_4_lut (.I0(n613), .I1(reset_per_frame_latched), .I2(write_to_dc32_fifo_latched_N_425), 
            .I3(n562[5]), .O(n2352));   // src/usb3_if.v(97[10] 190[8])
    defparam i1116_4_lut.LUT_INIT = 16'hcfdd;
    SB_LUT4 sub_113_add_2_3_lut (.I0(GND_net), .I1(num_lines_clocked_out[1]), 
            .I2(VCC_net), .I3(n10155), .O(num_lines_clocked_out_10__N_371[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_3 (.CI(n10155), .I0(num_lines_clocked_out[1]), 
            .I1(VCC_net), .CO(n10156));
    SB_LUT4 sub_113_add_2_2_lut (.I0(GND_net), .I1(num_lines_clocked_out[0]), 
            .I2(n1[0]), .I3(VCC_net), .O(num_lines_clocked_out_10__N_371[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_2 (.CI(VCC_net), .I0(num_lines_clocked_out[0]), 
            .I1(n1[0]), .CO(n10155));
    SB_LUT4 sub_113_add_2_12_lut (.I0(GND_net), .I1(num_lines_clocked_out[10]), 
            .I2(VCC_net), .I3(n10164), .O(num_lines_clocked_out_10__N_371[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_113_add_2_11_lut (.I0(GND_net), .I1(num_lines_clocked_out[9]), 
            .I2(VCC_net), .I3(n10163), .O(num_lines_clocked_out_10__N_371[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_11 (.CI(n10163), .I0(num_lines_clocked_out[9]), 
            .I1(VCC_net), .CO(n10164));
    SB_LUT4 sub_113_add_2_10_lut (.I0(GND_net), .I1(num_lines_clocked_out[8]), 
            .I2(VCC_net), .I3(n10162), .O(num_lines_clocked_out_10__N_371[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_10 (.CI(n10162), .I0(num_lines_clocked_out[8]), 
            .I1(VCC_net), .CO(n10163));
    SB_LUT4 sub_113_add_2_9_lut (.I0(GND_net), .I1(num_lines_clocked_out[7]), 
            .I2(VCC_net), .I3(n10161), .O(num_lines_clocked_out_10__N_371[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_9 (.CI(n10161), .I0(num_lines_clocked_out[7]), 
            .I1(VCC_net), .CO(n10162));
    SB_LUT4 sub_113_add_2_8_lut (.I0(GND_net), .I1(num_lines_clocked_out[6]), 
            .I2(VCC_net), .I3(n10160), .O(num_lines_clocked_out_10__N_371[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_8 (.CI(n10160), .I0(num_lines_clocked_out[6]), 
            .I1(VCC_net), .CO(n10161));
    SB_LUT4 sub_113_add_2_7_lut (.I0(GND_net), .I1(num_lines_clocked_out[5]), 
            .I2(VCC_net), .I3(n10159), .O(num_lines_clocked_out_10__N_371[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_7 (.CI(n10159), .I0(num_lines_clocked_out[5]), 
            .I1(VCC_net), .CO(n10160));
    SB_LUT4 sub_113_add_2_6_lut (.I0(GND_net), .I1(num_lines_clocked_out[4]), 
            .I2(VCC_net), .I3(n10158), .O(num_lines_clocked_out_10__N_371[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_6 (.CI(n10158), .I0(num_lines_clocked_out[4]), 
            .I1(VCC_net), .CO(n10159));
    SB_LUT4 sub_113_add_2_5_lut (.I0(GND_net), .I1(num_lines_clocked_out[3]), 
            .I2(VCC_net), .I3(n10157), .O(num_lines_clocked_out_10__N_371[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_5 (.CI(n10157), .I0(num_lines_clocked_out[3]), 
            .I1(VCC_net), .CO(n10158));
    SB_DFF state_FSM_i5 (.Q(n562[4]), .C(FIFO_CLK_c), .D(n4911));   // src/usb3_if.v(98[9] 189[16])
    SB_DFF state_FSM_i9 (.Q(n562[8]), .C(FIFO_CLK_c), .D(n4910));   // src/usb3_if.v(98[9] 189[16])
    SB_LUT4 sub_113_add_2_4_lut (.I0(GND_net), .I1(num_lines_clocked_out[2]), 
            .I2(VCC_net), .I3(n10156), .O(num_lines_clocked_out_10__N_371[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF dc32_fifo_data_in_latched__i1 (.Q(dc32_fifo_data_in_latched[0]), 
           .C(FIFO_CLK_c), .D(n4907));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i16 (.Q(dc32_fifo_data_in_latched[15]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D15_c_15), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i15 (.Q(dc32_fifo_data_in_latched[14]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D14_c_14), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i14 (.Q(dc32_fifo_data_in_latched[13]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D13_c_13), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i13 (.Q(dc32_fifo_data_in_latched[12]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D12_c_12), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i12 (.Q(dc32_fifo_data_in_latched[11]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D11_c_11), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i11 (.Q(dc32_fifo_data_in_latched[10]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D10_c_10), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i10 (.Q(dc32_fifo_data_in_latched[9]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D9_c_9), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i9 (.Q(dc32_fifo_data_in_latched[8]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D8_c_8), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i8 (.Q(dc32_fifo_data_in_latched[7]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D7_c_7), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i7 (.Q(dc32_fifo_data_in_latched[6]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D6_c_6), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i6 (.Q(dc32_fifo_data_in_latched[5]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D5_c_5), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i5 (.Q(dc32_fifo_data_in_latched[4]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D4_c_4), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i4 (.Q(dc32_fifo_data_in_latched[3]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D3_c_3), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i3 (.Q(dc32_fifo_data_in_latched[2]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D2_c_2), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i2 (.Q(dc32_fifo_data_in_latched[1]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D1_c_1), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_LUT4 i1_4_lut (.I0(n520), .I1(n562[1]), .I2(n562[0]), .I3(n551), 
            .O(n4));   // src/usb3_if.v(98[9] 189[16])
    defparam i1_4_lut.LUT_INIT = 16'heca0;
    SB_LUT4 i2_3_lut (.I0(n21), .I1(n4), .I2(n4224), .I3(GND_net), .O(n10282));   // src/usb3_if.v(98[9] 189[16])
    defparam i2_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i200_2_lut (.I0(dc32_fifo_almost_full), .I1(n562[5]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // src/usb3_if.v(98[9] 189[16])
    defparam i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1626_4_lut (.I0(n562[2]), .I1(n606), .I2(n524), .I3(dc32_fifo_empty_latched), 
            .O(n2992));   // src/usb3_if.v(98[9] 189[16])
    defparam i1626_4_lut.LUT_INIT = 16'hecee;
    SB_LUT4 i1635_4_lut (.I0(n562[6]), .I1(write_to_dc32_fifo_latched_N_425), 
            .I2(n551), .I3(n562[5]), .O(n3002));   // src/usb3_if.v(98[9] 189[16])
    defparam i1635_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 i212_2_lut (.I0(n551), .I1(n562[6]), .I2(GND_net), .I3(GND_net), 
            .O(n618));   // src/usb3_if.v(98[9] 189[16])
    defparam i212_2_lut.LUT_INIT = 16'h4444;
    SB_DFFN dc32_fifo_data_in_i16 (.Q(\dc32_fifo_data_in[15] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[15]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i15 (.Q(\dc32_fifo_data_in[14] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[14]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i14 (.Q(\dc32_fifo_data_in[13] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[13]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i13 (.Q(\dc32_fifo_data_in[12] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[12]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i12 (.Q(\dc32_fifo_data_in[11] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[11]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i11 (.Q(\dc32_fifo_data_in[10] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[10]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i10 (.Q(\dc32_fifo_data_in[9] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[9]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i9 (.Q(\dc32_fifo_data_in[8] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[8]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i8 (.Q(\dc32_fifo_data_in[7] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[7]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i7 (.Q(\dc32_fifo_data_in[6] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[6]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i6 (.Q(\dc32_fifo_data_in[5] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[5]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i5 (.Q(\dc32_fifo_data_in[4] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[4]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i4 (.Q(\dc32_fifo_data_in[3] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[3]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i3 (.Q(\dc32_fifo_data_in[2] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[2]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i2 (.Q(\dc32_fifo_data_in[1] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[1]));   // src/usb3_if.v(194[8] 197[4])
    SB_LUT4 i3_4_lut (.I0(state_timeout_counter[0]), .I1(state_timeout_counter[2]), 
            .I2(state_timeout_counter[1]), .I3(state_timeout_counter[3]), 
            .O(n524));   // src/usb3_if.v(151[21:49])
    defparam i3_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i2_3_lut_adj_1 (.I0(n524), .I1(n562[2]), .I2(dc32_fifo_empty_latched), 
            .I3(GND_net), .O(n4224));   // src/usb3_if.v(98[9] 189[16])
    defparam i2_3_lut_adj_1.LUT_INIT = 16'h4040;
    SB_DFFESR state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(FIFO_CLK_c), 
            .E(n4310), .D(n2400), .R(n4688));   // src/usb3_if.v(88[8] 191[4])
    SB_LUT4 i7_4_lut (.I0(num_lines_clocked_out[7]), .I1(num_lines_clocked_out[2]), 
            .I2(num_lines_clocked_out[9]), .I3(num_lines_clocked_out[0]), 
            .O(n18));   // src/usb3_if.v(175[29:57])
    defparam i7_4_lut.LUT_INIT = 16'hfeff;
    SB_DFFESS state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(FIFO_CLK_c), 
            .E(n4310), .D(n2401), .S(n4688));   // src/usb3_if.v(88[8] 191[4])
    SB_LUT4 i5_2_lut (.I0(num_lines_clocked_out[1]), .I1(num_lines_clocked_out[5]), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // src/usb3_if.v(175[29:57])
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut (.I0(num_lines_clocked_out[6]), .I1(n18), .I2(num_lines_clocked_out[3]), 
            .I3(num_lines_clocked_out[10]), .O(n20));   // src/usb3_if.v(175[29:57])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(FIFO_CLK_c), 
            .E(n4310), .D(n2402), .R(n4688));   // src/usb3_if.v(88[8] 191[4])
    SB_LUT4 i10_4_lut (.I0(num_lines_clocked_out[4]), .I1(n20), .I2(n16), 
            .I3(num_lines_clocked_out[8]), .O(n21));   // src/usb3_if.v(175[29:57])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1637_4_lut (.I0(n562[0]), .I1(n21), .I2(n522), .I3(n4224), 
            .O(n3004));   // src/usb3_if.v(98[9] 189[16])
    defparam i1637_4_lut.LUT_INIT = 16'hb3a0;
    SB_DFFSR write_to_dc32_fifo_latched_94 (.Q(write_to_dc32_fifo_latched), 
            .C(FIFO_CLK_c), .D(write_to_dc32_fifo_latched_N_425), .R(n2983));   // src/usb3_if.v(88[8] 191[4])
    SB_LUT4 i150_2_lut_3_lut (.I0(buffer_switch_done_latched), .I1(dc32_fifo_empty_latched), 
            .I2(DEBUG_1_c_c), .I3(GND_net), .O(n522));   // src/usb3_if.v(100[21:96])
    defparam i150_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i148_2_lut_3_lut (.I0(buffer_switch_done_latched), .I1(dc32_fifo_empty_latched), 
            .I2(DEBUG_1_c_c), .I3(GND_net), .O(n520));   // src/usb3_if.v(100[21:96])
    defparam i148_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i234_3_lut (.I0(n4181), .I1(FT_OE_N_420), .I2(n562[5]), .I3(GND_net), 
            .O(FT_OE_N_419));   // src/usb3_if.v(98[9] 189[16])
    defparam i234_3_lut.LUT_INIT = 16'hc5c5;
    SB_DFFESR num_lines_clocked_out_i1 (.Q(num_lines_clocked_out[1]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[1]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_LUT4 reduce_or_206_i1_2_lut (.I0(n562[8]), .I1(n562[4]), .I2(GND_net), 
            .I3(GND_net), .O(n613));   // src/usb3_if.v(98[9] 189[16])
    defparam reduce_or_206_i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i231_3_lut (.I0(n613), .I1(FT_OE_N_420), .I2(n562[5]), .I3(GND_net), 
            .O(FT_RD_N_422));   // src/usb3_if.v(98[9] 189[16])
    defparam i231_3_lut.LUT_INIT = 16'hc5c5;
    SB_DFFESR num_lines_clocked_out_i2 (.Q(num_lines_clocked_out[2]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[2]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR num_lines_clocked_out_i3 (.Q(num_lines_clocked_out[3]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[3]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR num_lines_clocked_out_i0 (.Q(num_lines_clocked_out[0]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[0]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR num_lines_clocked_out_i4 (.Q(num_lines_clocked_out[4]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[4]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR num_lines_clocked_out_i5 (.Q(num_lines_clocked_out[5]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[5]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_LUT4 sub_113_inv_0_i1_1_lut (.I0(dc32_fifo_empty_latched), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // src/usb3_if.v(174[50:77])
    defparam sub_113_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR num_lines_clocked_out_i6 (.Q(num_lines_clocked_out[6]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[6]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR num_lines_clocked_out_i7 (.Q(num_lines_clocked_out[7]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[7]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESS num_lines_clocked_out_i8 (.Q(num_lines_clocked_out[8]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[8]), .S(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR num_lines_clocked_out_i9 (.Q(num_lines_clocked_out[9]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[9]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESS num_lines_clocked_out_i10 (.Q(num_lines_clocked_out[10]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[10]), .S(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_CARRY sub_113_add_2_4 (.CI(n10156), .I0(num_lines_clocked_out[2]), 
            .I1(VCC_net), .CO(n10157));
    SB_DFFESR state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(FIFO_CLK_c), 
            .E(n4310), .D(n2399), .R(n4688));   // src/usb3_if.v(88[8] 191[4])
    SB_LUT4 i202_2_lut_3_lut_4_lut (.I0(n524), .I1(dc32_fifo_almost_full), 
            .I2(DEBUG_1_c_c), .I3(n562[1]), .O(n608));   // src/usb3_if.v(98[9] 189[16])
    defparam i202_2_lut_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1151_4_lut_4_lut (.I0(n562[5]), .I1(dc32_fifo_almost_full), 
            .I2(DEBUG_1_c_c), .I3(n524), .O(n2390));   // src/usb3_if.v(98[9] 189[16])
    defparam i1151_4_lut_4_lut.LUT_INIT = 16'h2276;
    SB_LUT4 i2_3_lut_4_lut (.I0(n575), .I1(n571), .I2(n562[8]), .I3(n562[4]), 
            .O(n4181));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1159_i2_4_lut (.I0(n2408), .I1(n3940), .I2(n2415), .I3(dc32_fifo_empty_latched), 
            .O(n2400));   // src/usb3_if.v(98[9] 189[16])
    defparam mux_1159_i2_4_lut.LUT_INIT = 16'h3f35;
    SB_LUT4 i1_2_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n3940));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10447_3_lut (.I0(n10783), .I1(reset_per_frame_latched), .I2(n4181), 
            .I3(GND_net), .O(n4310));   // src/usb3_if.v(97[10] 190[8])
    defparam i10447_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_4_lut_adj_2 (.I0(n562[0]), .I1(n2266), .I2(n520), .I3(DEBUG_1_c_c), 
            .O(n10783));   // src/usb3_if.v(97[10] 190[8])
    defparam i1_4_lut_adj_2.LUT_INIT = 16'h0ace;
    SB_LUT4 i3306_4_lut (.I0(n4310), .I1(n562[2]), .I2(n562[0]), .I3(n2390), 
            .O(n4688));   // src/usb3_if.v(88[8] 191[4])
    defparam i3306_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 i1050_2_lut (.I0(n562[5]), .I1(dc32_fifo_almost_full), .I2(GND_net), 
            .I3(GND_net), .O(n2266));
    defparam i1050_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_1159_i3_4_lut (.I0(n2408), .I1(n3938), .I2(n2415), .I3(n1[0]), 
            .O(n2401));   // src/usb3_if.v(98[9] 189[16])
    defparam mux_1159_i3_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 mux_1159_i4_4_lut (.I0(n12077), .I1(n3942), .I2(n2415), .I3(n2408), 
            .O(n2402));   // src/usb3_if.v(98[9] 189[16])
    defparam mux_1159_i4_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i10300_2_lut (.I0(n21), .I1(dc32_fifo_empty_latched), .I2(GND_net), 
            .I3(GND_net), .O(n12077));   // src/usb3_if.v(98[9] 189[16])
    defparam i10300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i179_2_lut_3_lut (.I0(n524), .I1(dc32_fifo_almost_full), .I2(DEBUG_1_c_c), 
            .I3(GND_net), .O(n551));   // src/usb3_if.v(155[26] 157[24])
    defparam i179_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1647_3_lut_4_lut (.I0(n562[5]), .I1(n562[8]), .I2(n562[4]), 
            .I3(FT_OE_N_420), .O(n3014));   // src/usb3_if.v(98[9] 189[16])
    defparam i1647_3_lut_4_lut.LUT_INIT = 16'hfcfe;
    SB_LUT4 i10389_2_lut (.I0(n562[5]), .I1(reset_per_frame_latched), .I2(GND_net), 
            .I3(GND_net), .O(n2983));   // src/usb3_if.v(88[8] 191[4])
    defparam i10389_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_3_lut (.I0(n524), .I1(reset_per_frame_latched), .I2(n562[2]), 
            .I3(GND_net), .O(n4486));
    defparam i1_3_lut.LUT_INIT = 16'hdcdc;
    SB_LUT4 mux_1159_i1_4_lut (.I0(n12030), .I1(state_timeout_counter[0]), 
            .I2(n2415), .I3(n2408), .O(n2399));   // src/usb3_if.v(98[9] 189[16])
    defparam mux_1159_i1_4_lut.LUT_INIT = 16'h3a3f;
    SB_LUT4 i10282_2_lut (.I0(n21), .I1(dc32_fifo_empty_latched), .I2(GND_net), 
            .I3(GND_net), .O(n12030));   // src/usb3_if.v(98[9] 189[16])
    defparam i10282_2_lut.LUT_INIT = 16'h4444;
    
endmodule

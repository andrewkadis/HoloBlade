// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Tue Sep 22 16:59:17 2020
//
// Verilog Description of module top
//

module top (ICE_SYSCLK, DCD, DSR, DTR, CTS, RST, UART_RX, UART_TX, 
            SEN, SCK, SOUT, SDAT, UPDATE, RESET, SLM_CLK, INVERT, 
            SYNC, VALID, DATA31, DATA0, DATA30, DATA29, DATA1, 
            DATA28, DATA27, DATA2, DATA26, DATA25, DATA3, DATA24, 
            DATA23, DATA4, DATA22, DATA21, DATA5, DATA20, DATA19, 
            DATA6, DATA18, DATA17, DATA7, DATA16, DATA15, DATA8, 
            DATA14, DATA13, DATA12, DATA11, DATA9, DATA10, FT_OE, 
            FT_RD, FT_WR, FT_SIWU, FR_RXF, FT_TXE, FIFO_BE3, FIFO_BE2, 
            FIFO_BE1, FIFO_BE0, FIFO_D31, FIFO_D30, FIFO_D29, FIFO_D28, 
            FIFO_D27, FIFO_CLK, FIFO_D26, FIFO_D25, FIFO_D24, FIFO_D23, 
            FIFO_D22, FIFO_D21, FIFO_D20, FIFO_D19, FIFO_D18, FIFO_D17, 
            FIFO_D16, FIFO_D15, FIFO_D14, FIFO_D13, FIFO_D12, FIFO_D11, 
            FIFO_D10, FIFO_D9, FIFO_D8, FIFO_D7, FIFO_D6, FIFO_D5, 
            FIFO_D4, FIFO_D3, FIFO_D2, FIFO_D1, FIFO_D0, DEBUG_0, 
            DEBUG_1, DEBUG_2, DEBUG_3, DEBUG_5, DEBUG_6, DEBUG_8, 
            DEBUG_9, ICE_CLK, ICE_CDONE, ICE_CREST) /* synthesis syn_module_defined=1 */ ;   // src/top.v(5[8:11])
    input ICE_SYSCLK;   // src/top.v(8[11:21])
    output DCD;   // src/top.v(11[12:15])
    output DSR;   // src/top.v(12[12:15])
    output DTR;   // src/top.v(13[12:15])
    output CTS;   // src/top.v(14[12:15])
    output RST;   // src/top.v(15[12:15])
    input UART_RX;   // src/top.v(16[12:19])
    output UART_TX;   // src/top.v(17[12:19])
    output SEN;   // src/top.v(20[12:15])
    output SCK;   // src/top.v(21[12:15])
    input SOUT;   // src/top.v(22[12:16])
    output SDAT;   // src/top.v(23[12:16])
    output UPDATE;   // src/top.v(27[12:18])
    output RESET;   // src/top.v(28[12:17])
    output SLM_CLK;   // src/top.v(29[12:19])
    output INVERT;   // src/top.v(30[12:18])
    output SYNC;   // src/top.v(31[12:16])
    output VALID;   // src/top.v(32[12:17])
    output DATA31;   // src/top.v(34[12:18])
    output DATA0;   // src/top.v(35[12:17])
    output DATA30;   // src/top.v(36[12:18])
    output DATA29;   // src/top.v(37[12:18])
    output DATA1;   // src/top.v(38[12:17])
    output DATA28;   // src/top.v(39[12:18])
    output DATA27;   // src/top.v(40[12:18])
    output DATA2;   // src/top.v(41[12:17])
    output DATA26;   // src/top.v(42[12:18])
    output DATA25;   // src/top.v(43[12:18])
    output DATA3;   // src/top.v(44[12:17])
    output DATA24;   // src/top.v(45[12:18])
    output DATA23;   // src/top.v(46[12:18])
    output DATA4;   // src/top.v(47[12:17])
    output DATA22;   // src/top.v(48[12:18])
    output DATA21;   // src/top.v(49[12:18])
    output DATA5;   // src/top.v(50[12:17])
    output DATA20;   // src/top.v(51[12:18])
    output DATA19;   // src/top.v(52[12:18])
    output DATA6;   // src/top.v(53[12:17])
    output DATA18;   // src/top.v(54[12:18])
    output DATA17;   // src/top.v(55[12:18])
    output DATA7;   // src/top.v(56[12:17])
    output DATA16;   // src/top.v(57[12:18])
    output DATA15;   // src/top.v(58[12:18])
    output DATA8;   // src/top.v(59[12:17])
    output DATA14;   // src/top.v(60[12:18])
    output DATA13;   // src/top.v(61[12:18])
    output DATA12;   // src/top.v(62[12:18])
    output DATA11;   // src/top.v(63[12:18])
    output DATA9;   // src/top.v(64[12:17])
    output DATA10;   // src/top.v(65[12:18])
    output FT_OE;   // src/top.v(69[12:17])
    output FT_RD;   // src/top.v(70[12:17])
    output FT_WR;   // src/top.v(71[12:17])
    output FT_SIWU;   // src/top.v(72[12:19])
    input FR_RXF;   // src/top.v(73[12:18])
    input FT_TXE;   // src/top.v(74[12:18])
    input FIFO_BE3;   // src/top.v(75[12:20])
    input FIFO_BE2;   // src/top.v(76[12:20])
    input FIFO_BE1;   // src/top.v(77[12:20])
    input FIFO_BE0;   // src/top.v(78[12:20])
    input FIFO_D31;   // src/top.v(79[12:20])
    input FIFO_D30;   // src/top.v(80[12:20])
    input FIFO_D29;   // src/top.v(81[12:20])
    input FIFO_D28;   // src/top.v(82[12:20])
    input FIFO_D27;   // src/top.v(83[12:20])
    input FIFO_CLK;   // src/top.v(84[12:20])
    input FIFO_D26;   // src/top.v(85[12:20])
    input FIFO_D25;   // src/top.v(86[12:20])
    input FIFO_D24;   // src/top.v(87[12:20])
    input FIFO_D23;   // src/top.v(88[12:20])
    input FIFO_D22;   // src/top.v(89[12:20])
    input FIFO_D21;   // src/top.v(90[12:20])
    input FIFO_D20;   // src/top.v(91[12:20])
    input FIFO_D19;   // src/top.v(92[12:20])
    input FIFO_D18;   // src/top.v(93[12:20])
    input FIFO_D17;   // src/top.v(94[12:20])
    input FIFO_D16;   // src/top.v(95[12:20])
    input FIFO_D15;   // src/top.v(97[11:19])
    input FIFO_D14;   // src/top.v(98[11:19])
    input FIFO_D13;   // src/top.v(99[11:19])
    input FIFO_D12;   // src/top.v(100[11:19])
    input FIFO_D11;   // src/top.v(101[11:19])
    input FIFO_D10;   // src/top.v(102[11:19])
    input FIFO_D9;   // src/top.v(103[11:18])
    input FIFO_D8;   // src/top.v(104[11:18])
    input FIFO_D7;   // src/top.v(105[11:18])
    input FIFO_D6;   // src/top.v(106[11:18])
    input FIFO_D5;   // src/top.v(107[11:18])
    input FIFO_D4;   // src/top.v(108[11:18])
    input FIFO_D3;   // src/top.v(109[11:18])
    input FIFO_D2;   // src/top.v(110[11:18])
    input FIFO_D1;   // src/top.v(111[11:18])
    input FIFO_D0;   // src/top.v(112[11:18])
    output DEBUG_0;   // src/top.v(115[12:19])
    output DEBUG_1;   // src/top.v(116[12:19])
    output DEBUG_2;   // src/top.v(117[12:19])
    output DEBUG_3;   // src/top.v(118[12:19])
    output DEBUG_5;   // src/top.v(119[12:19])
    output DEBUG_6;   // src/top.v(120[12:19])
    output DEBUG_8;   // src/top.v(121[12:19])
    output DEBUG_9;   // src/top.v(122[12:19])
    output ICE_CLK;   // src/top.v(125[12:19])
    output ICE_CDONE;   // src/top.v(126[12:21])
    output ICE_CREST;   // src/top.v(127[12:21])
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    
    wire GND_net, VCC_net, ICE_SYSCLK_c, UART_RX_c, UART_TX_c, SEN_c_1, 
<<<<<<< HEAD
        SCK_c_0, SOUT_c, SDAT_c_15, UPDATE_c_3, RESET_c, INVERT_c_4, 
        SYNC_c, VALID_c, FT_OE_c, FT_RD_c, FR_RXF_c, n11261, FIFO_D0_c_0, 
        DEBUG_0_c_24, DEBUG_1_c, DEBUG_3_c_0, DEBUG_5_c_0, DEBUG_6_c, 
        DEBUG_8_c, DEBUG_9_c, n11257, debug_led3, reset_all_w;
=======
<<<<<<< Updated upstream
        SCK_c_0, SOUT_c, SDAT_c_15, UPDATE_c_2, RESET_c, INVERT_c_3, 
        SYNC_c, DEBUG_9_c, DATA15_c, DEBUG_6_c, DATA14_c, DATA13_c, 
        DATA17_c, DATA12_c, DATA11_c, DATA18_c, DATA10_c, DATA9_c, 
        DATA19_c, DATA8_c, DATA7_c, DATA20_c, DATA6_c, DATA5_c, 
        FT_OE_c, DEBUG_2_c, DEBUG_1_c_c, FIFO_D15_c_15, FIFO_D14_c_14, 
        FIFO_D13_c_13, FIFO_D12_c_12, FIFO_D11_c_11, FIFO_D10_c_10, 
        FIFO_D9_c_9, FIFO_D8_c_8, FIFO_D7_c_7, FIFO_D6_c_6, FIFO_D5_c_5, 
        FIFO_D4_c_4, FIFO_D3_c_3, FIFO_D2_c_2, FIFO_D1_c_1, DEBUG_8_c_0_c, 
        DEBUG_0_c_24, DEBUG_3_c, DEBUG_5_c, debug_led3, reset_all_w;
>>>>>>> master
    wire [3:0]reset_clk_counter;   // src/top.v(242[10:27])
    
    wire reset_all, reset_per_frame, buffer_switch_done, dc32_fifo_full, 
        line_of_data_available, dc32_fifo_write_enable, dc32_fifo_read_enable, 
        sc32_fifo_read_enable;
    wire [3:0]state;   // src/timing_controller.v(78[11:16])
    
<<<<<<< HEAD
    wire n11239, sc32_fifo_almost_empty;
    wire [7:0]pc_data_rx;   // src/top.v(776[11:21])
=======
    wire dc32_fifo_almost_empty, get_next_word, \REG.mem_9_14 , \REG.mem_9_13 , 
        \REG.mem_9_12 , \REG.mem_9_11 , \REG.mem_9_10 , \REG.mem_9_9 , 
        \REG.mem_9_8 , \REG.mem_9_7 , \REG.mem_9_6 , \REG.mem_9_5 , 
        \REG.mem_9_4 , \REG.mem_9_3 , \REG.mem_9_2 , \REG.mem_9_1 , 
        \REG.mem_9_0 ;
    wire [31:0]fifo_data_out;   // src/top.v(545[12:25])
    wire [7:0]pc_data_rx;   // src/top.v(685[11:21])
=======
        SCK_c_0, SOUT_c, SDAT_c_15, UPDATE_c_3, RESET_c, INVERT_c_4, 
        SYNC_c, DEBUG_6_c, DATA31_c_31, DEBUG_8_c, DATA30_c_30, DATA29_c_29, 
        DATA1_c_1, DATA28_c_28, DATA27_c_27, DATA2_c_2, DATA26_c_26, 
        DATA25_c_25, DATA3_c_3, DATA24_c_24, DATA23_c_23, DATA4_c_4, 
        DATA22_c_22, DATA21_c_21, DATA5_c_5, DATA20_c_20, DATA19_c_19, 
        DATA6_c_6, DATA18_c_18, DATA17_c_17, DATA7_c_7, DATA16_c_16, 
        DATA15_c_15, DATA8_c_8, DATA14_c_14, DATA13_c_13, DATA12_c_12, 
        DATA11_c_11, DATA9_c_9, DATA10_c_10, FT_OE_c, FT_RD_c, FR_RXF_c, 
        FIFO_D31_c_31, FIFO_D30_c_30, FIFO_D29_c_29, FIFO_D28_c_28, 
        FIFO_D27_c_27, FIFO_D26_c_26, FIFO_D25_c_25, FIFO_D24_c_24, 
        FIFO_D23_c_23, FIFO_D22_c_22, FIFO_D21_c_21, FIFO_D20_c_20, 
        FIFO_D19_c_19, FIFO_D18_c_18, FIFO_D17_c_17, FIFO_D16_c_16, 
        FIFO_D15_c_15, FIFO_D14_c_14, FIFO_D13_c_13, FIFO_D12_c_12, 
        FIFO_D11_c_11, FIFO_D10_c_10, FIFO_D9_c_9, FIFO_D8_c_8, FIFO_D7_c_7, 
        FIFO_D6_c_6, FIFO_D5_c_5, FIFO_D4_c_4, FIFO_D3_c_3, FIFO_D2_c_2, 
        FIFO_D1_c_1, DEBUG_3_c_0_c, DEBUG_0_c_24, DEBUG_1_c, DEBUG_2_c, 
        DEBUG_5_c_0, DEBUG_9_c_0, debug_led3, n8, reset_all_w;
    wire [3:0]reset_clk_counter;   // src/top.v(242[10:27])
    
    wire reset_all, reset_per_frame, buffer_switch_done, dc32_fifo_full, 
        line_of_data_available, dc32_fifo_write_enable;
    wire [31:0]dc32_fifo_data_in;   // src/top.v(541[13:30])
    
    wire dc32_fifo_empty, dc32_fifo_almost_empty, dc32_fifo_read_enable;
    wire [31:0]dc32_fifo_data_out;   // src/top.v(483[23:41])
    
    wire sc32_fifo_read_enable;
    wire [3:0]state;   // src/timing_controller.v(78[11:16])
    
    wire sc32_fifo_almost_empty;
    wire [7:0]pc_data_rx;   // src/top.v(776[11:21])
>>>>>>> Stashed changes
>>>>>>> master
    
    wire tx_uart_active_flag, spi_start_transfer_r, multi_byte_spi_trans_flag_r;
    wire [7:0]tx_addr_byte;   // src/top.v(898[11:23])
    wire [7:0]tx_data_byte;   // src/top.v(900[11:23])
    wire [7:0]rx_buf_byte;   // src/top.v(907[11:22])
    
    wire is_tx_fifo_full_flag, fifo_write_cmd, spi_rx_byte_ready, fifo_read_cmd, 
        is_fifo_empty_flag;
    wire [31:0]fifo_temp_output;   // src/top.v(997[12:28])
    
    wire even_byte_flag, uart_rx_complete_rising_edge, uart_rx_complete_prev, 
<<<<<<< HEAD
        reset_all_w_N_61, n5734, start_tx_N_64, pll_clk_unbuf, multi_byte_spi_trans_flag_r_N_72, 
        \REG.mem_13_0 , \REG.mem_1_0 , \REG.mem_22_0 , \REG.mem_21_0 , 
        \REG.mem_20_0 , \REG.mem_19_0 , \REG.mem_18_0 , \REG.mem_12_0 , 
        n5731, n5730, buffer_switch_done_latched, \REG.mem_15_0 , n1967, 
        \REG.mem_24_0 , n1459, n11193, n59, n47, n10373, n5726, 
        n5725, n5724, n5723, n5721, n5720, n5719, n5718, n5717, 
        n5716, n5715, n5714, n5713, n5712, \REG.mem_5_0 , \REG.mem_11_0 ;
    wire [7:0]state_timeout_counter_adj_1430;   // src/bluejay_data.v(52[11:32])
=======
<<<<<<< Updated upstream
        \REG.mem_15_14 , reset_all_w_N_61, \REG.mem_11_8 , \REG.mem_11_7 , 
        start_tx_N_64, pll_clk_unbuf, n7386;
    wire [3:0]state;   // src/timing_controller.v(51[11:16])
>>>>>>> master
    
    wire n80, n10372, n10371, n5711, n5710, n5709, n5708, n5707, 
        n5706, n5705, n5704, n5703, n5702, n5701, n5700, n5699, 
        n5698, n5697, n5696, n5695, n2329, n5694, n5693, n5692, 
        n5691, n5690, n5689, n5688, n5687, n5686, n5685, n5684, 
        bluejay_data_out_31__N_919, bluejay_data_out_31__N_920, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // src/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // src/uart_rx.v(36[17:26])
    
    wire n5683, n5682, n5681, n5679, n5677, n5675, n5674, n10370, 
        n5673, n5672, n5671, n5670, n5669, n5668, n5667;
    wire [2:0]r_SM_Main_2__N_949;
    
    wire n5666, n5665, n10369, n18, n25;
    wire [2:0]r_SM_Main_adj_1435;   // src/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_1437;   // src/uart_tx.v(33[16:27])
    wire [7:0]r_Tx_Data;   // src/uart_tx.v(34[16:25])
    wire [2:0]r_SM_Main_2__N_1028;
    wire [2:0]r_SM_Main_2__N_1025;
    
    wire n106, n24, n5664, n5663, n5662, n5661, \REG.mem_14_0 , 
        n10368;
    wire [15:0]tx_shift_reg;   // src/spi.v(70[12:24])
    wire [15:0]rx_shift_reg;   // src/spi.v(72[12:24])
    
    wire n11094, n10367, n10366, n10365, n10364, n5659, n10209, 
        n10363, n2072, n5658, n5657, n5656, n10362, n11171, n10361, 
        n10360, n10359, n5655, n5654, n5653, n5652, n5651, n5650, 
        n5649, n5648, n10358, n5132, n10357, \REG.mem_10_0 , n10356, 
        n2704, \REG.mem_16_0 , n11046, \REG.mem_9_0 ;
    wire [5:0]wr_addr_r;   // src/fifo_dc_32_lut_gen.v(196[29:38])
    wire [5:0]wr_addr_nxt_c;   // src/fifo_dc_32_lut_gen.v(198[29:42])
    wire [5:0]rp_sync1_r;   // src/fifo_dc_32_lut_gen.v(201[37:47])
    wire [5:0]wr_grey_w;   // src/fifo_dc_32_lut_gen.v(203[38:47])
    wire [5:0]wr_grey_sync_r;   // src/fifo_dc_32_lut_gen.v(204[37:51])
    wire [5:0]rd_addr_r;   // src/fifo_dc_32_lut_gen.v(217[29:38])
    wire [5:0]rd_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(221[30:42])
    wire [5:0]wp_sync1_r;   // src/fifo_dc_32_lut_gen.v(222[37:47])
    wire [5:0]rd_grey_sync_r;   // src/fifo_dc_32_lut_gen.v(225[37:51])
    
    wire n5645, rd_fifo_en_w, \aempty_flag_impl.ae_flag_nxt_w , \REG.mem_4_0 , 
        n10355, n11079, n10354;
    wire [5:0]rd_addr_nxt_c_5__N_572;
    
    wire n5644, n5643, \REG.mem_8_0 , n5120, n10353, n63, n5113, 
        n10352, n10351, \REG.mem_7_0 , n5504, wr_fifo_en_w, rd_fifo_en_prev_r;
    wire [2:0]wr_addr_r_adj_1490;   // src/fifo_quad_word_mod.v(65[31:40])
    wire [2:0]wr_addr_p1_w_adj_1492;   // src/fifo_quad_word_mod.v(67[32:44])
    wire [2:0]rd_addr_r_adj_1493;   // src/fifo_quad_word_mod.v(69[31:40])
    wire [2:0]rd_addr_p1_w_adj_1495;   // src/fifo_quad_word_mod.v(71[32:44])
    
    wire \REG.mem_3_0 , n10350;
    wire [31:0]\mem_LUT.data_raw_r ;   // src/fifo_quad_word_mod.v(449[42:52])
    
    wire n32, empty_o_N_1333, n3254, n15, n5101, \REG.mem_6_0 , 
        n10640, \REG.mem_2_0 , n3426, n24_adj_1400, n5081, n11863, 
        n5642, n5641, n5640, \REG.mem_17_0 , \REG.mem_0_0 , n5639, 
        n5500, \REG.mem_23_0 , \REG.mem_25_0 , \REG.mem_26_0 , \REG.mem_27_0 , 
        \REG.mem_28_0 , \REG.mem_29_0 , n8057, n11700, \REG.mem_30_0 , 
        n6690, \REG.mem_31_0 , n10668, n7, n6, n5638, n23, n5637, 
        n5214, n5212, n5019, n5457, n5527, n7836, n5825, n10381, 
        n11101, n5821, n11362, n3, n5817, n25_adj_1401, n11691, 
        n8012, n5812, n5808, n5635, n5634, n5633, n5632, n5631, 
        n5628, n5626, n5625, n5624, n5623, n5622, n5621, n5620, 
        n5618, n5617, n5616, n5615, n5614, n5611, n5610, n5607, 
        n5525, n21, n30, n22, n31, n23_adj_1402, n32_adj_1403, 
        n24_adj_1404, n33, n25_adj_1405, n34, n26, n35, n27, n28, 
        n29, n4, n20, n5159, n130, n129, n128, n127, n126, 
        n125, n124, n123, n122, n121, n120, n119, n118, n117, 
        n116, n115, n114, n113, n112, n111, n110, n109, n108, 
        n107, n106_adj_1406, n5605, n5769, n5766, n5762, n5761, 
        n5758, n5757, n5756, n5755, n5752, n5751, n5750, n5749, 
        n5748, n5745, n5742, n5741, n5738, n5735, n10792, n4_adj_1407, 
        n6_adj_1408, n5, n13, n2, n22_adj_1409, n23_adj_1410, n11, 
        n10, n3_adj_1411, n10608, n4943, n7_adj_1412, n4715, n16, 
        n17, n10471, n4_adj_1413, n10469, n21_adj_1414, n9, n12, 
        n4_adj_1415, n20_adj_1416, n14, n15_adj_1417, n4_adj_1418, 
        n10467, n1, n19, n8;
    
    VCC i2 (.Y(VCC_net));
    timing_controller timing_controller_inst (.SLM_CLK_c(SLM_CLK_c), .GND_net(GND_net), 
            .sc32_fifo_read_enable(sc32_fifo_read_enable), .n10668(n10668), 
            .VCC_net(VCC_net), .state({state}), .dc32_fifo_read_enable(dc32_fifo_read_enable), 
            .n1967(n1967), .DEBUG_8_c(DEBUG_8_c), .DEBUG_6_c(DEBUG_6_c), 
            .n63(n63), .n5132(n5132), .\state_timeout_counter[7] (state_timeout_counter_adj_1430[7]), 
            .n3(n3), .n11094(n11094), .n5500(n5500), .n1459(n1459), 
            .n106(n106), .n80(n80), .n5504(n5504), .buffer_switch_done(buffer_switch_done), 
            .n2072(n2072), .n7836(n7836), .INVERT_c_4(INVERT_c_4), .n11257(n11257), 
            .dc32_fifo_full(dc32_fifo_full), .n11101(n11101), .n7(n7), 
            .n59(n59), .n6(n6), .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .n4943(n4943), .n47(n47), .reset_all(reset_all), .n11700(n11700), 
            .reset_per_frame(reset_per_frame), .n8057(n8057), .line_of_data_available(line_of_data_available), 
            .UPDATE_c_3(UPDATE_c_3)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(472[19] 493[2])
    SB_DFF uart_rx_complete_prev_83 (.Q(uart_rx_complete_prev), .C(SLM_CLK_c), 
<<<<<<< HEAD
           .D(debug_led3));   // src/top.v(1156[8] 1162[4])
    SB_LUT4 i4242_3_lut (.I0(rx_shift_reg[6]), .I1(rx_shift_reg[5]), .I2(n5113), 
            .I3(GND_net), .O(n5701));   // src/spi.v(76[8] 221[4])
    defparam i4242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(is_fifo_empty_flag), .I1(fifo_write_cmd), .I2(n32), 
            .I3(GND_net), .O(n24_adj_1400));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i4243_3_lut (.I0(rx_shift_reg[5]), .I1(rx_shift_reg[4]), .I2(n5113), 
            .I3(GND_net), .O(n5702));   // src/spi.v(76[8] 221[4])
    defparam i4243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9595_4_lut (.I0(rd_addr_p1_w_adj_1495[2]), .I1(n11863), .I2(wr_addr_r_adj_1490[2]), 
            .I3(wr_addr_r_adj_1490[1]), .O(n11171));
    defparam i9595_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i4244_3_lut (.I0(rx_shift_reg[4]), .I1(rx_shift_reg[3]), .I2(n5113), 
            .I3(GND_net), .O(n5703));   // src/spi.v(76[8] 221[4])
    defparam i4244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4245_3_lut (.I0(rx_shift_reg[3]), .I1(rx_shift_reg[2]), .I2(n5113), 
            .I3(GND_net), .O(n5704));   // src/spi.v(76[8] 221[4])
    defparam i4245_3_lut.LUT_INIT = 16'hcaca;
    bluejay_data bluejay_data_inst (.VCC_net(VCC_net), .VALID_c(VALID_c), 
            .SLM_CLK_c(SLM_CLK_c), .bluejay_data_out_31__N_920(bluejay_data_out_31__N_920), 
            .buffer_switch_done(buffer_switch_done), .GND_net(GND_net), 
            .n1459(n1459), .n3(n3), .buffer_switch_done_latched(buffer_switch_done_latched), 
            .n5132(n5132), .n80(n80), .n11094(n11094), .SYNC_c(SYNC_c), 
            .bluejay_data_out_31__N_919(bluejay_data_out_31__N_919), .\state_timeout_counter[7] (state_timeout_counter_adj_1430[7]), 
            .line_of_data_available(line_of_data_available), .n5504(n5504), 
            .n5500(n5500), .sc32_fifo_almost_empty(sc32_fifo_almost_empty), 
            .n5616(n5616), .DEBUG_8_c(DEBUG_8_c), .n106(n106)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(717[14] 730[2])
    SB_GB clk_gb (.GLOBAL_BUFFER_OUTPUT(SLM_CLK_c), .USER_SIGNAL_TO_GLOBAL_BUFFER(pll_clk_unbuf)) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=222, LSE_RLINE=228 */ ;   // src/clock.v(82[7:96])
=======
           .D(debug_led3));   // src/top.v(1065[8] 1071[4])
    bluejay_data bluejay_data_inst (.dc32_fifo_almost_full(dc32_fifo_almost_full), 
            .n771(n771), .dc32_fifo_almost_empty(dc32_fifo_almost_empty), 
            .bluejay_data_out_31__N_736(bluejay_data_out_31__N_736), .buffer_switch_done_latched(buffer_switch_done_latched), 
            .GND_net(GND_net), .DEBUG_9_c(DEBUG_9_c), .SLM_CLK_c(SLM_CLK_c), 
            .DATA19_c(DATA19_c), .buffer_switch_done(buffer_switch_done), 
            .n4937(n4937), .DATA18_c(DATA18_c), .n4936(n4936), .DATA17_c(DATA17_c), 
            .n6112(n6112), .DEBUG_6_c(DEBUG_6_c), .DATA15_c(DATA15_c), 
            .DATA14_c(DATA14_c), .DATA13_c(DATA13_c), .DATA12_c(DATA12_c), 
            .n843(n843), .VCC_net(VCC_net), .DATA11_c(DATA11_c), .DATA10_c(DATA10_c), 
            .SYNC_c(SYNC_c), .bluejay_data_out_31__N_737(bluejay_data_out_31__N_737), 
            .n10277(n10277), .DATA9_c(DATA9_c), .DATA8_c(DATA8_c), .DATA7_c(DATA7_c), 
            .DATA6_c(DATA6_c), .\rd_sig_diff0_w[1] (rd_sig_diff0_w[1]), 
            .get_next_word(get_next_word), .\rd_sig_diff0_w[0] (rd_sig_diff0_w[0]), 
            .\rd_sig_diff0_w[2] (rd_sig_diff0_w[2]), .n10873(n10873), .n10877(n10877), 
            .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .DATA5_c(DATA5_c), .DATA20_c(DATA20_c), .\fifo_data_out[4] (fifo_data_out[4]), 
            .\fifo_data_out[5] (fifo_data_out[5]), .\fifo_data_out[6] (fifo_data_out[6]), 
            .\fifo_data_out[7] (fifo_data_out[7]), .\fifo_data_out[11] (fifo_data_out[11]), 
            .\fifo_data_out[10] (fifo_data_out[10]), .\fifo_data_out[3] (fifo_data_out[3]), 
            .\fifo_data_out[15] (fifo_data_out[15]), .\fifo_data_out[14] (fifo_data_out[14]), 
            .\fifo_data_out[13] (fifo_data_out[13]), .\fifo_data_out[12] (fifo_data_out[12]), 
            .\fifo_data_out[9] (fifo_data_out[9]), .\fifo_data_out[8] (fifo_data_out[8])) /* synthesis syn_module_defined=1 */ ;   // src/top.v(626[14] 639[2])
    SB_LUT4 i4128_3_lut (.I0(\REG.mem_36_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n29), .I3(GND_net), .O(n5511));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4128_3_lut.LUT_INIT = 16'hcaca;
    SB_GB clk_gb (.GLOBAL_BUFFER_OUTPUT(SLM_CLK_c), .USER_SIGNAL_TO_GLOBAL_BUFFER(pll_clk_unbuf)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=222, LSE_RLINE=228 */ ;   // src/clock.v(82[7:96])
    SB_LUT4 i4129_3_lut (.I0(\REG.mem_36_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n29), .I3(GND_net), .O(n5512));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4130_3_lut (.I0(\REG.mem_36_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n29), .I3(GND_net), .O(n5513));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4131_3_lut (.I0(\REG.mem_36_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n29), .I3(GND_net), .O(n5514));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4131_3_lut.LUT_INIT = 16'hcaca;
=======
        get_next_word, reset_all_w_N_61, n13008, start_tx_N_64, pll_clk_unbuf, 
        multi_byte_spi_trans_flag_r_N_72, \REG.mem_11_16 , \REG.mem_11_15 , 
        \REG.mem_11_14 , \REG.mem_11_13 , \REG.mem_11_12 , \REG.mem_11_11 , 
        \REG.mem_11_10 , \REG.mem_11_9 , \REG.mem_11_8 , \REG.mem_11_7 , 
        \REG.mem_11_6 , \REG.mem_11_5 , \REG.mem_11_4 , \REG.mem_11_3 , 
        \REG.mem_11_2 , \REG.mem_11_1 , \REG.mem_22_6 , \REG.mem_22_5 , 
        \REG.mem_20_29 , \REG.mem_20_28 , \REG.mem_20_27 , \REG.mem_20_26 , 
        \REG.mem_20_25 , \REG.mem_20_24 , \REG.mem_20_23 , \REG.mem_20_22 , 
        \REG.mem_20_21 , \REG.mem_20_20 , \REG.mem_20_19 , \REG.mem_20_18 , 
        \REG.mem_20_17 , n5343, \REG.mem_20_16 , \REG.mem_20_15 , \REG.mem_20_14 , 
        \REG.mem_20_13 , \REG.mem_20_12 , \REG.mem_20_11 , \REG.mem_20_10 , 
        \REG.mem_20_9 , \REG.mem_20_8 , \REG.mem_20_7 , \REG.mem_20_6 , 
        \REG.mem_20_5 , \REG.mem_11_0 , \REG.mem_10_31 , \REG.mem_10_30 , 
        \REG.mem_10_29 , \REG.mem_10_28 , \REG.mem_10_27 , \REG.mem_20_4 , 
        \REG.mem_20_3 , \REG.mem_20_2 , \REG.mem_20_1 , \REG.mem_20_0 , 
        \REG.mem_17_31 , \REG.mem_17_30 , \REG.mem_17_29 , \REG.mem_17_28 , 
        \REG.mem_17_27 , \REG.mem_17_26 , \REG.mem_17_25 , \REG.mem_17_24 , 
        \REG.mem_17_23 , \REG.mem_17_22 , \REG.mem_17_21 , \REG.mem_17_20 , 
        \REG.mem_17_19 , \REG.mem_17_18 , \REG.mem_17_17 , \REG.mem_17_16 , 
        \REG.mem_17_15 , \REG.mem_17_14 , \REG.mem_17_13 , \REG.mem_17_12 , 
        \REG.mem_17_11 , \REG.mem_17_10 , \REG.mem_17_9 , \REG.mem_17_8 , 
        \REG.mem_17_7 , \REG.mem_17_6 , \REG.mem_17_5 , \REG.mem_17_4 , 
        \REG.mem_17_3 , \REG.mem_17_2 , \REG.mem_17_1 , \REG.mem_17_0 , 
        \REG.mem_10_26 , \REG.mem_10_25 , \REG.mem_10_24 , \REG.mem_10_23 , 
        \REG.mem_10_22 , \REG.mem_10_21 , \REG.mem_10_20 , \REG.mem_10_19 , 
        \REG.mem_10_18 , \REG.mem_10_17 , \REG.mem_10_16 , \REG.mem_10_15 , 
        \REG.mem_10_14 , \REG.mem_10_13 , \REG.mem_10_12 , \REG.mem_10_11 , 
        \REG.mem_10_10 , \REG.mem_10_9 , \REG.mem_10_8 , \REG.mem_10_7 , 
        \REG.mem_10_6 , \REG.mem_10_5 , \REG.mem_10_4 , \REG.mem_10_3 , 
        \REG.mem_10_2 , \REG.mem_10_1 , \REG.mem_10_0 , \REG.mem_9_31 , 
        \REG.mem_9_30 , \REG.mem_9_29 , \REG.mem_9_28 , \REG.mem_9_27 , 
        reset_per_frame_latched, buffer_switch_done_latched, n2407, \REG.mem_22_4 , 
        \REG.mem_22_3 , \REG.mem_22_2 , n12261, n2335, \REG.mem_22_1 , 
        \REG.mem_22_0 , \REG.mem_21_31 , \REG.mem_21_30 , n5366, \REG.mem_21_29 , 
        \REG.mem_21_28 , n5365, n5350, n2075, \REG.mem_21_27 , \REG.mem_21_26 , 
        \REG.mem_21_25 , n5665, n5662, n5659, n5656, n5653, \REG.mem_9_26 , 
        \REG.mem_9_25 , \REG.mem_9_24 , \REG.mem_9_23 , \REG.mem_9_22 , 
        \REG.mem_4_25 , \REG.mem_4_24 , \REG.mem_4_23 , \REG.mem_4_22 , 
        \REG.mem_4_21 , \REG.mem_4_20 , \REG.mem_4_19 , \REG.mem_4_18 , 
        \REG.mem_4_17 , \REG.mem_4_16 , \REG.mem_4_15 , \REG.mem_4_14 , 
        \REG.mem_4_13 , \REG.mem_4_12 , \REG.mem_4_11 , \REG.mem_4_10 , 
        \REG.mem_4_9 , \REG.mem_4_8 , \REG.mem_4_7 , \REG.mem_4_6 , 
        \REG.mem_4_5 , \REG.mem_4_4 , \REG.mem_4_3 , \REG.mem_4_2 , 
        \REG.mem_4_1 , \REG.mem_4_0 , \REG.mem_21_24 , \REG.mem_21_23 , 
        \REG.mem_21_22 , \REG.mem_21_21 , n5338, n5344, n5346, n5354, 
        n5356, n5364, n5648, n5645, n5636, n5635, \REG.mem_9_21 , 
        \REG.mem_9_20 , \REG.mem_9_19 , \REG.mem_9_18 , \REG.mem_9_17 , 
        \REG.mem_9_16 , \REG.mem_9_15 , \REG.mem_9_14 , bluejay_data_out_31__N_920, 
        bluejay_data_out_31__N_921, bluejay_data_out_31__N_922, \REG.mem_21_20 , 
        r_Rx_Data;
    wire [2:0]r_Bit_Index;   // src/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main_adj_1467;   // src/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_1469;   // src/uart_tx.v(33[16:27])
    wire [7:0]r_Tx_Data;   // src/uart_tx.v(34[16:25])
    wire [2:0]r_SM_Main_2__N_1029;
    wire [2:0]r_SM_Main_2__N_1026;
    
    wire n12978;
    wire [15:0]tx_shift_reg;   // src/spi.v(70[12:24])
    wire [15:0]rx_shift_reg;   // src/spi.v(72[12:24])
    
    wire n4688, n2180, \REG.mem_11_31 , n5615, n5611, n5086, \REG.mem_9_13 , 
        \REG.mem_9_12 , \REG.mem_9_11 , \REG.mem_9_10 , \REG.mem_9_9 , 
        \REG.mem_9_8 , \REG.mem_9_7 , \REG.mem_9_6 , \REG.mem_9_5 , 
        \REG.mem_9_4 , \REG.mem_9_3 , \REG.mem_9_2 , \REG.mem_9_1 , 
        \REG.mem_9_0 , \REG.mem_8_31 , \REG.mem_8_30 , n5610, \REG.mem_21_19 , 
        \REG.mem_21_18 , \REG.mem_11_30 , n5608, n5607, \REG.mem_11_29 , 
        \REG.mem_11_28 , \REG.mem_11_27 , \REG.mem_11_26 , \REG.mem_11_25 , 
        \REG.mem_11_24 , n5604, \REG.mem_11_23 , \REG.mem_11_22 , \REG.mem_11_21 , 
        \REG.mem_11_20 , n5603, n5602, \REG.mem_21_17 , n5337, \REG.mem_8_29 , 
        \REG.mem_8_28 , \REG.mem_8_27 , \REG.mem_8_26 , \REG.mem_8_25 , 
        \REG.mem_8_24 , \REG.mem_8_23 , \REG.mem_8_22 , \REG.mem_8_21 , 
        \REG.mem_8_20 , \REG.mem_8_19 , \REG.mem_8_18 , \REG.mem_8_17 , 
        \REG.mem_8_16 , \REG.mem_8_15 , \REG.mem_8_14 , \REG.mem_8_13 , 
        \REG.mem_8_12 , \REG.mem_8_11 , \REG.mem_8_10 , \REG.mem_8_9 , 
        \REG.mem_8_8 , \REG.mem_8_7 , \REG.mem_8_6 ;
    wire [5:0]wr_addr_r;   // src/fifo_dc_32_lut_gen.v(196[29:38])
    wire [5:0]wr_addr_nxt_c;   // src/fifo_dc_32_lut_gen.v(198[29:42])
    wire [5:0]wr_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(200[30:42])
    wire [5:0]rp_sync1_r;   // src/fifo_dc_32_lut_gen.v(201[37:47])
    wire [5:0]wr_grey_sync_r;   // src/fifo_dc_32_lut_gen.v(204[37:51])
    
    wire \REG.mem_11_19 , \REG.mem_11_18 , \REG.mem_11_17 ;
    wire [5:0]wp_sync1_r;   // src/fifo_dc_32_lut_gen.v(222[37:47])
    wire [5:0]rd_grey_sync_r;   // src/fifo_dc_32_lut_gen.v(225[37:51])
    
    wire wr_fifo_en_w, \aempty_flag_impl.ae_flag_nxt_w , n5600;
    wire [5:0]rd_addr_nxt_c_5__N_573;
    
    wire \REG.mem_8_5 , \REG.mem_8_4 , \REG.mem_8_3 , \REG.mem_8_2 , 
        \REG.mem_8_1 , \REG.mem_8_0 , \REG.mem_7_31 , \REG.mem_7_30 , 
        \REG.mem_7_29 , \REG.mem_7_28 , \REG.mem_7_27 , \REG.mem_7_26 , 
        \REG.mem_7_25 , \REG.mem_7_24 , \REG.mem_7_23 , \REG.mem_7_22 , 
        \REG.mem_7_21 , \REG.mem_7_20 , \REG.mem_7_19 , \REG.mem_7_18 , 
        \REG.mem_7_17 , \REG.mem_7_16 , \REG.mem_7_15 , \REG.mem_7_14 , 
        \REG.mem_7_13 , \REG.mem_7_12 , \REG.mem_7_11 , \REG.mem_7_10 , 
        \REG.mem_7_9 , \REG.mem_7_8 , \REG.mem_7_7 , \REG.mem_7_6 , 
        \REG.mem_21_16 , \REG.mem_21_15 , n663, \REG.mem_7_5 , \REG.mem_7_4 , 
        \REG.mem_7_3 , \REG.mem_7_2 , \REG.mem_7_1 , \REG.mem_7_0 , 
        \REG.mem_6_31 , \REG.mem_6_30 , \REG.mem_6_29 , \REG.mem_6_28 , 
        \REG.mem_6_27 , \REG.mem_6_26 , \REG.mem_6_25 , \REG.mem_6_24 , 
        \REG.mem_6_23 , \REG.mem_6_22 , \REG.mem_6_21 , \REG.mem_6_20 , 
        \REG.mem_6_19 , \REG.mem_6_18 , \REG.mem_6_17 , \REG.mem_6_16 , 
        \REG.mem_6_15 , \REG.mem_6_14 , \REG.mem_6_13 , \REG.mem_6_12 , 
        \REG.mem_6_11 , \REG.mem_6_10 , \REG.mem_6_9 , \REG.mem_6_8 , 
        \REG.mem_6_7 , \REG.mem_6_6 , wr_fifo_en_w_adj_1416, rd_fifo_en_w, 
        rd_fifo_en_prev_r;
    wire [2:0]wr_addr_r_adj_1517;   // src/fifo_quad_word_mod.v(65[31:40])
    wire [2:0]wr_addr_p1_w_adj_1519;   // src/fifo_quad_word_mod.v(67[32:44])
    wire [2:0]rd_addr_r_adj_1520;   // src/fifo_quad_word_mod.v(69[31:40])
    wire [2:0]rd_addr_p1_w_adj_1522;   // src/fifo_quad_word_mod.v(71[32:44])
    wire [31:0]\mem_LUT.data_raw_r ;   // src/fifo_quad_word_mod.v(449[42:52])
    
    wire \REG.mem_6_5 , \REG.mem_6_4 , \REG.mem_6_3 , \REG.mem_6_2 , 
        \REG.mem_6_1 , \REG.mem_6_0 , n5599, n3353, \REG.mem_5_31 , 
        \REG.mem_5_30 , \REG.mem_5_29 , \REG.mem_5_28 , \REG.mem_5_27 , 
        \REG.mem_5_26 , \REG.mem_5_25 , \REG.mem_5_24 , \REG.mem_5_23 , 
        \REG.mem_5_22 , \REG.mem_5_21 , \REG.mem_5_20 , \REG.mem_5_19 , 
        \REG.mem_5_18 , \REG.mem_5_17 , \REG.mem_5_16 , \REG.mem_5_15 , 
        \REG.mem_5_14 , \REG.mem_5_13 , \REG.mem_5_12 , \REG.mem_5_11 , 
        \REG.mem_5_10 , \REG.mem_5_9 , \REG.mem_5_8 , \REG.mem_5_7 , 
        \REG.mem_5_6 , \REG.mem_5_5 , \REG.mem_5_4 , \REG.mem_5_3 , 
        \REG.mem_5_2 , \REG.mem_5_1 , \REG.mem_5_0 , \REG.mem_1_31 , 
        \REG.mem_1_30 , \REG.mem_1_29 , \REG.mem_1_28 , \REG.mem_1_27 , 
        \REG.mem_1_26 , \REG.mem_1_25 , \REG.mem_1_24 , \REG.mem_1_23 , 
        \REG.mem_1_22 , \REG.mem_1_21 , \REG.mem_1_20 , \REG.mem_1_19 , 
        \REG.mem_1_18 , \REG.mem_1_17 , \REG.mem_1_16 , \REG.mem_1_15 , 
        \REG.mem_1_14 , \REG.mem_1_13 , \REG.mem_1_12 , \REG.mem_1_11 , 
        \REG.mem_1_10 , \REG.mem_1_9 , \REG.mem_1_8 , \REG.mem_1_7 , 
        \REG.mem_1_6 , \REG.mem_1_5 , \REG.mem_1_4 , \REG.mem_4_31 , 
        \REG.mem_4_30 , \REG.mem_4_29 , \REG.mem_4_28 , \REG.mem_4_27 , 
        \REG.mem_4_26 , n3468, \REG.mem_1_3 , \REG.mem_1_2 , \REG.mem_1_1 , 
        \REG.mem_1_0 , n8_adj_1418, n5596, n5595, n5594, n5593, 
        n934, n5592, n5590, n5589, n5339, n1013, \REG.mem_21_14 , 
        n5347, n12177, \REG.mem_21_13 , \REG.mem_21_12 , n5348, \REG.mem_21_11 , 
        n5367, \REG.mem_21_10 , \REG.mem_21_9 , \REG.mem_21_8 , \REG.mem_21_7 , 
        \REG.mem_21_6 , \REG.mem_21_5 , \REG.mem_21_4 , \REG.mem_21_3 , 
        \REG.mem_21_2 , \REG.mem_21_1 , \REG.mem_21_0 , \REG.mem_20_31 , 
        n5588, \REG.mem_20_30 , n5587, n5586, n12882, \REG.mem_22_7 , 
        \REG.mem_22_8 , \REG.mem_22_9 , \REG.mem_22_10 , \REG.mem_22_11 , 
        \REG.mem_22_12 , \REG.mem_22_13 , \REG.mem_22_14 , \REG.mem_22_15 , 
        \REG.mem_22_16 , \REG.mem_22_17 , \REG.mem_22_18 , \REG.mem_22_19 , 
        \REG.mem_22_20 , \REG.mem_22_21 , \REG.mem_22_22 , \REG.mem_22_23 , 
        \REG.mem_22_24 , \REG.mem_22_25 , \REG.mem_22_26 , \REG.mem_22_27 , 
        \REG.mem_22_28 , \REG.mem_22_29 , \REG.mem_22_30 , \REG.mem_22_31 , 
        \REG.mem_23_0 , \REG.mem_23_1 , \REG.mem_23_2 , \REG.mem_23_3 , 
        \REG.mem_23_4 , \REG.mem_23_5 , \REG.mem_23_6 , \REG.mem_23_7 , 
        \REG.mem_23_8 , \REG.mem_23_9 , \REG.mem_23_10 , \REG.mem_23_11 , 
        \REG.mem_23_12 , \REG.mem_23_13 , \REG.mem_23_14 , \REG.mem_23_15 , 
        \REG.mem_23_16 , \REG.mem_23_17 , \REG.mem_23_18 , \REG.mem_23_19 , 
        \REG.mem_23_20 , \REG.mem_23_21 , \REG.mem_23_22 , \REG.mem_23_23 , 
        \REG.mem_23_24 , \REG.mem_23_25 , \REG.mem_23_26 , \REG.mem_23_27 , 
        \REG.mem_23_28 , \REG.mem_23_29 , \REG.mem_23_30 , \REG.mem_23_31 , 
        \REG.mem_24_0 , \REG.mem_24_1 , \REG.mem_24_2 , \REG.mem_24_3 , 
        \REG.mem_24_4 , \REG.mem_24_5 , \REG.mem_24_6 , \REG.mem_24_7 , 
        \REG.mem_24_8 , \REG.mem_24_9 , \REG.mem_24_10 , \REG.mem_24_11 , 
        \REG.mem_24_12 , \REG.mem_24_13 , \REG.mem_24_14 , \REG.mem_24_15 , 
        \REG.mem_24_16 , \REG.mem_24_17 , \REG.mem_24_18 , \REG.mem_24_19 , 
        \REG.mem_24_20 , \REG.mem_24_21 , \REG.mem_24_22 , \REG.mem_24_23 , 
        \REG.mem_24_24 , \REG.mem_24_25 , \REG.mem_24_26 , \REG.mem_24_27 , 
        \REG.mem_24_28 , \REG.mem_24_29 , \REG.mem_24_30 , \REG.mem_24_31 , 
        \REG.mem_25_0 , \REG.mem_25_1 , \REG.mem_25_2 , \REG.mem_25_3 , 
        \REG.mem_25_4 , \REG.mem_25_5 , \REG.mem_25_6 , \REG.mem_25_7 , 
        \REG.mem_25_8 , \REG.mem_25_9 , \REG.mem_25_10 , \REG.mem_25_11 , 
        \REG.mem_25_12 , \REG.mem_25_13 , \REG.mem_25_14 , \REG.mem_25_15 , 
        \REG.mem_25_16 , \REG.mem_25_17 , \REG.mem_25_18 , \REG.mem_25_19 , 
        \REG.mem_25_20 , \REG.mem_25_21 , \REG.mem_25_22 , \REG.mem_25_23 , 
        \REG.mem_25_24 , \REG.mem_25_25 , \REG.mem_25_26 , \REG.mem_25_27 , 
        \REG.mem_25_28 , \REG.mem_25_29 , \REG.mem_25_30 , \REG.mem_25_31 , 
        \REG.mem_26_0 , \REG.mem_26_1 , \REG.mem_26_2 , \REG.mem_26_3 , 
        \REG.mem_26_4 , \REG.mem_26_5 , \REG.mem_26_6 , \REG.mem_26_7 , 
        \REG.mem_26_8 , \REG.mem_26_9 , \REG.mem_26_10 , \REG.mem_26_11 , 
        \REG.mem_26_12 , \REG.mem_26_13 , \REG.mem_26_14 , \REG.mem_26_15 , 
        \REG.mem_26_16 , \REG.mem_26_17 , \REG.mem_26_18 , \REG.mem_26_19 , 
        \REG.mem_26_20 , \REG.mem_26_21 , \REG.mem_26_22 , \REG.mem_26_23 , 
        \REG.mem_26_24 , \REG.mem_26_25 , \REG.mem_26_26 , \REG.mem_26_27 , 
        \REG.mem_26_28 , \REG.mem_26_29 , \REG.mem_26_30 , \REG.mem_26_31 , 
        \REG.mem_27_0 , \REG.mem_27_1 , \REG.mem_27_2 , \REG.mem_27_3 , 
        \REG.mem_27_4 , \REG.mem_27_5 , \REG.mem_27_6 , \REG.mem_27_7 , 
        \REG.mem_27_8 , \REG.mem_27_9 , \REG.mem_27_10 , \REG.mem_27_11 , 
        \REG.mem_27_12 , \REG.mem_27_13 , \REG.mem_27_14 , \REG.mem_27_15 , 
        \REG.mem_27_16 , \REG.mem_27_17 , \REG.mem_27_18 , \REG.mem_27_19 , 
        \REG.mem_27_20 , \REG.mem_27_21 , \REG.mem_27_22 , \REG.mem_27_23 , 
        \REG.mem_27_24 , \REG.mem_27_25 , \REG.mem_27_26 , \REG.mem_27_27 , 
        \REG.mem_27_28 , \REG.mem_27_29 , \REG.mem_27_30 , \REG.mem_27_31 , 
        n6, n7, n8_adj_1419, n9, n10, n11, n12, n13, n16, 
        n22, n23, n24, n25, n26, n27, n28, n29, n32, n9015, 
        n9013, n12176, n12175, n15, n12477, n12439, n7_adj_1420, 
        n12836, n7021, n7020, n7019, n7018, n7017, n7016, n7015, 
        n7014, n7013, n7012, n7011, n7010, n7009, n7008, n7007, 
        n7006, n7005, n7004, n7003, n7002, n7000, n6998, n6997, 
        n6996, n6995, n6994, n6993, n6992, n6991, n6990, n6989, 
        n6988, n6987, n6986, n6985, n6984, n6983, n6982, n6981, 
        n6980, n6979, n6978, n6977, n6976, n6975, n6968, n6967, 
        n6966, n6965, n6964, n6963, n6962, n6961, n6960, n6956, 
        n13052, n6950, n6947, n6941, n6938, n6937, n6936, n6935, 
        n6934, n6933, n6932, n6930, n6928, n6923, n6920, n6909, 
        n6908, n6907, n6906, n6905, n6904, n6903, n6493, n6492, 
        n6491, n6490, n6489, n6488, n6487, n6486, n6485, n6484, 
        n6483, n6482, n6481, n6480, n6479, n6478, n6477, n6476, 
        n6475, n6474, n6473, n6472, n6471, n6470, n6469, n6468, 
        n6467, n6466, n6465, n6464, n6463, n6462, n6461, n6460, 
        n6459, n6458, n6457, n6456, n6455, n6454, n6453, n6452, 
        n6451, n6450, n6449, n6448, n6447, n6446, n6445, n6444, 
        n6443, n6442, n6441, n6440, n6439, n6438, n6437, n6436, 
        n6435, n6434, n6433, n6432, n6431, n6430, n6429, n6428, 
        n6427, n6426, n6425, n6424, n6423, n6422, n6421, n6420, 
        n6419, n6418, n6417, n6416, n6415, n6414, n6413, n6412, 
        n6411, n6410, n6409, n6408, n6407, n6406, n6405, n6404, 
        n6403, n6402, n6401, n6400, n6399, n6398, n6397, n6396, 
        n6395, n6394, n6393, n6392, n6391, n6390, n6389, n6388, 
        n6387, n6386, n6385, n6384, n6383, n6382, n6381, n6380, 
        n6379, n6378, n6377, n6376, n6375, n6374, n6373, n6372, 
        n6371, n6370, n6369, n6368, n6367, n6366, n6365, n6364, 
        n6363, n6362, n6361, n6360, n6359, n6358, n6357, n6356, 
        n6355, n6354, n6353, n6352, n6351, n6350, n6349, n6348, 
        n6347, n6346, n6345, n6344, n6343, n6342, n6341, n6340, 
        n6339, n6338, n6337, n6336, n6335, n6334, n6333, n6332, 
        n6331, n6330, n6329, n6328, n6327, n6326, n6325, n6324, 
        n6323, n6322, n6321, n6320, n6319, n6318, n6317, n6316, 
        n6315, n6314, n6313, n6312, n6311, n6310, n6309, n6308, 
        n6307, n6306, n6305, n6304, n6303, n6302, n6301, n6300, 
        n6299, n6298, n6297, n6296, n6295, n6294, n6293, n6292, 
        n6291, n6290, n6289, n6288, n6287, n6286, n6285, n6284, 
        n6283, n6282, n6281, n6280, n6279, n6278, n6277, n6276, 
        n6275, n6274, n6273, n6272, n6271, n6270, n6269, n6268, 
        n6267, n6266, n6265, n6264, n6263, n6262, n6261, n6260, 
        n6259, n6258, n6257, n6256, n6255, n6254, n6253, n6252, 
        n6251, n6250, n6249, n6248, n6247, n6246, n6245, n6244, 
        n6243, n6242, n6241, n6240, n6239, n6238, n6173, n6172, 
        n6171, n6170, n6169, n6168, n6167, n6166, n6165, n6164, 
        n6163, n6162, n6161, n6160, n6159, n6158, n6157, n6156, 
        n6155, n6154, n6153, n6152, n6151, n6150, n6149, n6148, 
        n6147, n6146, n6145, n6144, n6143, n6142, n5981, n5980, 
        n5979, n5978, n5977, n5976, n5975, n5974, n5973, n5972, 
        n5971, n5970, n5969, n5968, n5967, n5966, n5965, n5964, 
        n5963, n5962, n5961, n5960, n5959, n5958, n5957, n5956, 
        n5955, n5954, n5953, n5952, n5951, n5950, n5949, n5948, 
        n5947, n5946, n5945, n5944, n5943, n5942, n5941, n5940, 
        n5939, n5938, n5937, n5936, n5935, n5934, n5933, n5932, 
        n5931, n5930, n5929, n5928, n5927, n5926, n5925, n5924, 
        n5923, n5922, n5921, n5920, n5919, n5918, n5917, n5916, 
        n5915, n5914, n5362, n5024, n130, n129, n128, n127, 
        n126, n125, n124, n123, n122, n121, n120, n119, n118, 
        n117, n5913, n5912, n5911, n5910, n5909, n5908, n5907, 
        n5906, n24_adj_1421, n23_adj_1422, n22_adj_1423, n21, n20, 
        n19, n18, n17, n16_adj_1424, n15_adj_1425, n14, n13_adj_1426, 
        n12_adj_1427, n11_adj_1428, n10_adj_1429, n9_adj_1430, n8_adj_1431, 
        n7_adj_1432, n6_adj_1433, n5, n4, n3, n2, n5905, n5904, 
        n5903, n5902, n5901, n5900, n5899, n5898, n63, n5360, 
        n5897, n5896, n5460, n5895, n5894, n5893, n5892, n5891, 
        n5890, n5889, n5888, n5887, n5886, n5885, n5884, n5883, 
        n5882, n5881, n5880, n5879, n5878, n5877, n5876, n5875, 
        n5874, n5873, n5872, n5871, n5870, n5869, n5868, n5867, 
        n5866, n5865, n5864, n5863, n5862, n5861, n5860, n5859, 
        n5858, n5857, n5856, n5855, n5854, n5853, n5852, n5851, 
        n116, n115, n5850, n114, n113, n112, n5849, n107, n5848, 
        n5847, n106, n111, n110, n109, n108, n5846, n5845, n5844, 
        n5843, n5842, n5841, n5840, n5839, n5838, n5837, n5836, 
        n5341, n5835, n5834, n5833, n5832, n5342, n5831, n5830, 
        n5358, n5829, n5828, n5827, n5357, n5826, n5825, n5824, 
        n5823, n5822, n5821, n5820, n5819, n5818, n5817, n5816, 
        n5815, n5814, n5813, n5812, n5811, n5810, n5809, n5808, 
        n5807, n5806, n5805, n5804, n5803, n5802, n5801, n5800, 
        n5799, n5798, n5797, n4_adj_1434, n5796, n5795, n5794, 
        n5793, n5792, n5791, n5790, n5789, n5788, n5787, n5786, 
        n5785, n5784, n5783, n5782, n5781, n5780, n5779, n5778, 
        n5777, n5776, n5775, n4903, n5774, n5345, n5773, n5772, 
        n5771, n5770, n5769, n5768, n4_adj_1435, n5767, n5766, 
        n5765, n5764, n5763, n5762, n4_adj_1436, n5761, n5760, 
        n5759, n5758, n5757, n5756, n5755, n5754, n5753, n5752, 
        n5751, n5750, n5749, n5748, n5747, n5746, n5745, n25_adj_1437, 
        n5744, n5743, n4884, n5585, n5583, n5582, n5581, n5580, 
        n5578, n5577, n5576, n5742, n5741, n5740, n5739, n5738, 
        n5737, n5736, n5735, n5734, n5733, n5575, n5574, n5573, 
        n5572, n5571, n5567, n5732, n5731, n5730, n5729, n5728, 
        n5727, n5726, n5363, n12174, n12173, n5565, n5564, n5560, 
        n5559, n5558, n5557, n5556, n25_adj_1438, n5361, n12215, 
        n5359, n12172, n12171, n12170, n12169, n12168, n12167, 
        n12166, n12165, n12164, n12163, n12162, n12161, n12160, 
        n5384, n8_adj_1439, n12159, n12158, n5555, n5353, n12157, 
        n12156, n12155, n12154, n5554, n5352, n3963, n5355, n12964, 
        n12040, n12938, n12906, n14242, n32_adj_1440, n4_adj_1441, 
        n4_adj_1442, n13034, n5340, n5349, n24_adj_1443, n5552, 
        n5551, n5550, n4794, n8659, n5351, n4837, n4314, n25_adj_1444, 
        n12884, n4790, n12310, n4787, n12308, n12537, n12304, 
        n4446, n16231;
    
    VCC i2 (.Y(VCC_net));
    timing_controller timing_controller_inst (.SLM_CLK_c(SLM_CLK_c), .DEBUG_2_c(DEBUG_2_c), 
            .sc32_fifo_read_enable(sc32_fifo_read_enable), .state({state}), 
            .dc32_fifo_read_enable(dc32_fifo_read_enable), .n63(n63), .GND_net(GND_net), 
            .VCC_net(VCC_net), .n2075(n2075), .n2180(n2180), .n9015(n9015), 
            .buffer_switch_done(buffer_switch_done), .n12477(n12477), .n8659(n8659), 
            .reset_all(reset_all), .line_of_data_available(line_of_data_available), 
            .n7(n7_adj_1420), .n8(n8_adj_1439), .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .INVERT_c_4(INVERT_c_4), .n4903(n4903), .get_next_word(get_next_word), 
            .dc32_fifo_almost_empty(dc32_fifo_almost_empty), .n4688(n4688), 
            .dc32_fifo_full(dc32_fifo_full), .n9013(n9013), .n12884(n12884), 
            .reset_per_frame(reset_per_frame), .UPDATE_c_3(UPDATE_c_3), 
            .n25(n25_adj_1444), .n12882(n12882)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(472[19] 493[2])
    SB_LUT4 i4974_3_lut (.I0(\REG.mem_26_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n7), .I3(GND_net), .O(n6448));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5486_3_lut (.I0(r_Tx_Data[1]), .I1(fifo_temp_output[1]), .I2(n4314), 
            .I3(GND_net), .O(n6960));   // src/uart_tx.v(38[10] 141[8])
    defparam i5486_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF fifo_read_cmd_80 (.Q(fifo_read_cmd), .C(SLM_CLK_c), .D(start_tx_N_64));   // src/top.v(1001[8] 1019[4])
    bluejay_data bluejay_data_inst (.VCC_net(VCC_net), .DEBUG_6_c(DEBUG_6_c), 
            .SLM_CLK_c(SLM_CLK_c), .GND_net(GND_net), .n4903(n4903), .buffer_switch_done(buffer_switch_done), 
            .n6968(n6968), .DEBUG_8_c(DEBUG_8_c), .buffer_switch_done_latched(buffer_switch_done_latched), 
            .n934(n934), .n12261(n12261), .n1013(n1013), .bluejay_data_out_31__N_920(bluejay_data_out_31__N_920), 
            .bluejay_data_out_31__N_921(bluejay_data_out_31__N_921), .bluejay_data_out_31__N_922(bluejay_data_out_31__N_922), 
            .SYNC_c(SYNC_c), .DATA10_c_10(DATA10_c_10), .n5367(n5367), 
            .line_of_data_available(line_of_data_available), .DATA9_c_9(DATA9_c_9), 
            .n5366(n5366), .DATA11_c_11(DATA11_c_11), .n5365(n5365), .DATA12_c_12(DATA12_c_12), 
            .n5364(n5364), .DATA13_c_13(DATA13_c_13), .n5363(n5363), .DATA14_c_14(DATA14_c_14), 
            .n5362(n5362), .DATA8_c_8(DATA8_c_8), .n5361(n5361), .DATA15_c_15(DATA15_c_15), 
            .n5360(n5360), .DATA16_c_16(DATA16_c_16), .n5359(n5359), .DATA7_c_7(DATA7_c_7), 
            .n5358(n5358), .DATA17_c_17(DATA17_c_17), .n5357(n5357), .DATA18_c_18(DATA18_c_18), 
            .n5356(n5356), .DATA6_c_6(DATA6_c_6), .n5355(n5355), .DATA19_c_19(DATA19_c_19), 
            .n5354(n5354), .DATA20_c_20(DATA20_c_20), .n5353(n5353), .DATA5_c_5(DATA5_c_5), 
            .n5352(n5352), .DATA21_c_21(DATA21_c_21), .n5351(n5351), .DATA22_c_22(DATA22_c_22), 
            .n5350(n5350), .DATA4_c_4(DATA4_c_4), .n5349(n5349), .DATA23_c_23(DATA23_c_23), 
            .n5348(n5348), .DATA24_c_24(DATA24_c_24), .n5347(n5347), .DATA3_c_3(DATA3_c_3), 
            .n5346(n5346), .DATA25_c_25(DATA25_c_25), .n5345(n5345), .DATA26_c_26(DATA26_c_26), 
            .n5344(n5344), .DATA2_c_2(DATA2_c_2), .n5343(n5343), .DATA27_c_27(DATA27_c_27), 
            .n5342(n5342), .n5573(n5573), .get_next_word(get_next_word), 
            .DATA28_c_28(DATA28_c_28), .n5341(n5341), .DATA1_c_1(DATA1_c_1), 
            .n5340(n5340), .DATA29_c_29(DATA29_c_29), .n5339(n5339), .DATA30_c_30(DATA30_c_30), 
            .n5338(n5338), .DATA31_c_31(DATA31_c_31), .n5337(n5337), .sc32_fifo_almost_empty(sc32_fifo_almost_empty)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(717[14] 730[2])
    SB_LUT4 i4975_3_lut (.I0(\REG.mem_26_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n7), .I3(GND_net), .O(n6449));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4975_3_lut.LUT_INIT = 16'hcaca;
    SB_GB clk_gb (.GLOBAL_BUFFER_OUTPUT(SLM_CLK_c), .USER_SIGNAL_TO_GLOBAL_BUFFER(pll_clk_unbuf)) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=222, LSE_RLINE=228 */ ;   // src/clock.v(82[7:96])
    SB_LUT4 i4976_3_lut (.I0(\REG.mem_26_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n7), .I3(GND_net), .O(n6450));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4976_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF uart_rx_complete_prev_83 (.Q(uart_rx_complete_prev), .C(SLM_CLK_c), 
           .D(debug_led3));   // src/top.v(1156[8] 1162[4])
>>>>>>> Stashed changes
>>>>>>> master
    SB_IO RST_pad (.PACKAGE_PIN(RST), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RST_pad.PIN_TYPE = 6'b011001;
    defparam RST_pad.PULLUP = 1'b0;
    defparam RST_pad.NEG_TRIGGER = 1'b0;
    defparam RST_pad.IO_STANDARD = "SB_LVCMOS";
<<<<<<< HEAD
    SB_LUT4 i4246_3_lut (.I0(rx_shift_reg[2]), .I1(rx_shift_reg[1]), .I2(n5113), 
            .I3(GND_net), .O(n5705));   // src/spi.v(76[8] 221[4])
    defparam i4246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4247_3_lut (.I0(rx_shift_reg[1]), .I1(rx_shift_reg[0]), .I2(n5113), 
            .I3(GND_net), .O(n5706));   // src/spi.v(76[8] 221[4])
    defparam i4247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(reset_all_w), .I1(n11171), .I2(n24_adj_1400), 
            .I3(n4), .O(n11046));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut.LUT_INIT = 16'hfbfa;
    SB_LUT4 i4248_4_lut (.I0(\REG.mem_19_0 ), .I1(DEBUG_3_c_0), .I2(n27), 
            .I3(wr_addr_r[4]), .O(n5707));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4248_4_lut.LUT_INIT = 16'hcaaa;
    SB_DFF tx_data_byte_r_i0_i1 (.Q(tx_data_byte[1]), .C(SLM_CLK_c), .D(n5730));   // src/top.v(1165[8] 1232[4])
    SB_LUT4 i4169_3_lut (.I0(tx_addr_byte[0]), .I1(tx_data_byte[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5628));   // src/top.v(1165[8] 1232[4])
    defparam i4169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4249_4_lut (.I0(\REG.mem_20_0 ), .I1(DEBUG_3_c_0), .I2(n29), 
            .I3(wr_addr_r[4]), .O(n5708));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4249_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i4172_4_lut (.I0(\REG.mem_1_0 ), .I1(DEBUG_3_c_0), .I2(n23_adj_1402), 
            .I3(wr_addr_r[4]), .O(n5631));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4172_4_lut.LUT_INIT = 16'haaca;
=======
<<<<<<< Updated upstream
    SB_LUT4 i3515_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4898));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i3515_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4624_3_lut (.I0(\REG.mem_63_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n2), .I3(GND_net), .O(n6007));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4625_3_lut (.I0(\REG.mem_63_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n2), .I3(GND_net), .O(n6008));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4132_3_lut (.I0(\REG.mem_36_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n29), .I3(GND_net), .O(n5515));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4133_3_lut (.I0(\REG.mem_36_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n29), .I3(GND_net), .O(n5516));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4134_3_lut (.I0(\REG.mem_36_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n29), .I3(GND_net), .O(n5517));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4135_3_lut (.I0(\REG.mem_36_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n29), .I3(GND_net), .O(n5518));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4626_3_lut (.I0(\REG.mem_63_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n2), .I3(GND_net), .O(n6009));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4627_3_lut (.I0(\REG.mem_63_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n2), .I3(GND_net), .O(n6010));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4136_3_lut (.I0(\REG.mem_36_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n29), .I3(GND_net), .O(n5519));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4137_3_lut (.I0(\REG.mem_36_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n29), .I3(GND_net), .O(n5520));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4198_3_lut (.I0(\REG.mem_39_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n26), .I3(GND_net), .O(n5581));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4138_3_lut (.I0(\REG.mem_36_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n29), .I3(GND_net), .O(n5521));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4139_3_lut (.I0(\REG.mem_36_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n29), .I3(GND_net), .O(n5522));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4199_3_lut (.I0(\REG.mem_39_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n26), .I3(GND_net), .O(n5582));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4140_3_lut (.I0(\REG.mem_36_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n29), .I3(GND_net), .O(n5523));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4141_3_lut (.I0(\REG.mem_36_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n29), .I3(GND_net), .O(n5524));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4141_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_all_r_77 (.Q(reset_all_w), .C(SLM_CLK_c), .D(reset_all_w_N_61));   // src/top.v(246[8] 264[4])
    SB_LUT4 i4200_3_lut (.I0(\REG.mem_39_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n26), .I3(GND_net), .O(n5583));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4142_3_lut (.I0(\REG.mem_36_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n29), .I3(GND_net), .O(n5525));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4143_3_lut (.I0(\REG.mem_36_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n29), .I3(GND_net), .O(n5526));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4144_3_lut (.I0(tx_addr_byte[7]), .I1(tx_data_byte[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5527));   // src/top.v(1074[8] 1141[4])
    defparam i4144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4201_3_lut (.I0(\REG.mem_39_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n26), .I3(GND_net), .O(n5584));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4145_3_lut (.I0(tx_addr_byte[6]), .I1(tx_data_byte[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5528));   // src/top.v(1074[8] 1141[4])
    defparam i4145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4628_3_lut (.I0(\REG.mem_63_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n2), .I3(GND_net), .O(n6011));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4202_3_lut (.I0(\REG.mem_39_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n26), .I3(GND_net), .O(n5585));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4146_3_lut (.I0(tx_addr_byte[5]), .I1(tx_data_byte[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5529));   // src/top.v(1074[8] 1141[4])
    defparam i4146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4203_3_lut (.I0(\REG.mem_39_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n26), .I3(GND_net), .O(n5586));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4147_3_lut (.I0(tx_addr_byte[4]), .I1(tx_data_byte[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5530));   // src/top.v(1074[8] 1141[4])
    defparam i4147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4148_3_lut (.I0(tx_addr_byte[3]), .I1(tx_data_byte[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5531));   // src/top.v(1074[8] 1141[4])
    defparam i4148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4149_3_lut (.I0(tx_addr_byte[2]), .I1(tx_data_byte[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5532));   // src/top.v(1074[8] 1141[4])
    defparam i4149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4204_3_lut (.I0(\REG.mem_39_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n26), .I3(GND_net), .O(n5587));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4205_3_lut (.I0(\REG.mem_39_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n26), .I3(GND_net), .O(n5588));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4629_3_lut (.I0(\REG.mem_63_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n2), .I3(GND_net), .O(n6012));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4630_3_lut (.I0(\REG.mem_63_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n2), .I3(GND_net), .O(n6013));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4631_3_lut (.I0(\REG.mem_63_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n2), .I3(GND_net), .O(n6014));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4150_3_lut (.I0(tx_addr_byte[1]), .I1(tx_data_byte[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5533));   // src/top.v(1074[8] 1141[4])
    defparam i4150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4157_3_lut (.I0(\REG.mem_37_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n28), .I3(GND_net), .O(n5540));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4632_3_lut (.I0(\REG.mem_63_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n2), .I3(GND_net), .O(n6015));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4158_3_lut (.I0(\REG.mem_37_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n28), .I3(GND_net), .O(n5541));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4159_3_lut (.I0(\REG.mem_37_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n28), .I3(GND_net), .O(n5542));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4160_3_lut (.I0(\REG.mem_37_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n28), .I3(GND_net), .O(n5543));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4161_3_lut (.I0(\REG.mem_37_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n28), .I3(GND_net), .O(n5544));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4162_3_lut (.I0(\REG.mem_37_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n28), .I3(GND_net), .O(n5545));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4163_3_lut (.I0(\REG.mem_37_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n28), .I3(GND_net), .O(n5546));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4164_3_lut (.I0(\REG.mem_37_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n28), .I3(GND_net), .O(n5547));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4165_3_lut (.I0(\REG.mem_37_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n28), .I3(GND_net), .O(n5548));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4633_3_lut (.I0(\REG.mem_63_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n2), .I3(GND_net), .O(n6016));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4206_3_lut (.I0(\REG.mem_39_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n26), .I3(GND_net), .O(n5589));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [13]), .I3(fifo_data_out[13]), .O(n10580));
    defparam i12_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4634_3_lut (.I0(\REG.mem_63_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n2), .I3(GND_net), .O(n6017));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4166_3_lut (.I0(\REG.mem_37_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n28), .I3(GND_net), .O(n5549));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4167_3_lut (.I0(\REG.mem_37_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n28), .I3(GND_net), .O(n5550));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4168_3_lut (.I0(\REG.mem_37_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n28), .I3(GND_net), .O(n5551));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4278_3_lut (.I0(\REG.mem_44_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n21), .I3(GND_net), .O(n5661));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4207_3_lut (.I0(\REG.mem_40_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n25), .I3(GND_net), .O(n5590));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4169_3_lut (.I0(\REG.mem_37_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n28), .I3(GND_net), .O(n5552));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4279_3_lut (.I0(\REG.mem_44_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n21), .I3(GND_net), .O(n5662));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4170_3_lut (.I0(\REG.mem_37_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n28), .I3(GND_net), .O(n5553));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4171_3_lut (.I0(\REG.mem_37_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n28), .I3(GND_net), .O(n5554));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4208_3_lut (.I0(\REG.mem_40_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n25), .I3(GND_net), .O(n5591));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4172_3_lut (.I0(\REG.mem_37_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n28), .I3(GND_net), .O(n5555));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4173_3_lut (.I0(\REG.mem_38_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n27), .I3(GND_net), .O(n5556));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4175_3_lut (.I0(\REG.mem_38_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n27), .I3(GND_net), .O(n5558));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4176_3_lut (.I0(\REG.mem_38_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n27), .I3(GND_net), .O(n5559));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4177_3_lut (.I0(\REG.mem_38_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n27), .I3(GND_net), .O(n5560));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_74 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [14]), .I3(fifo_data_out[14]), .O(n10582));
    defparam i12_4_lut_4_lut_adj_74.LUT_INIT = 16'h3120;
    SB_LUT4 i4178_3_lut (.I0(\REG.mem_38_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n27), .I3(GND_net), .O(n5561));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4179_3_lut (.I0(\REG.mem_38_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n27), .I3(GND_net), .O(n5562));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4180_3_lut (.I0(\REG.mem_38_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n27), .I3(GND_net), .O(n5563));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4181_3_lut (.I0(\REG.mem_38_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n27), .I3(GND_net), .O(n5564));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4182_3_lut (.I0(\REG.mem_38_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n27), .I3(GND_net), .O(n5565));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4183_3_lut (.I0(\REG.mem_38_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n27), .I3(GND_net), .O(n5566));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4184_3_lut (.I0(\REG.mem_38_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n27), .I3(GND_net), .O(n5567));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4209_3_lut (.I0(\REG.mem_40_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n25), .I3(GND_net), .O(n5592));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4185_3_lut (.I0(\REG.mem_38_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n27), .I3(GND_net), .O(n5568));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4186_3_lut (.I0(\REG.mem_38_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n27), .I3(GND_net), .O(n5569));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4281_3_lut (.I0(\REG.mem_44_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n21), .I3(GND_net), .O(n5664));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4282_3_lut (.I0(\REG.mem_44_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n21), .I3(GND_net), .O(n5665));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4210_3_lut (.I0(\REG.mem_40_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n25), .I3(GND_net), .O(n5593));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4187_3_lut (.I0(\REG.mem_38_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n27), .I3(GND_net), .O(n5570));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4211_3_lut (.I0(\REG.mem_40_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n25), .I3(GND_net), .O(n5594));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4212_3_lut (.I0(\REG.mem_40_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n25), .I3(GND_net), .O(n5595));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4188_3_lut (.I0(\REG.mem_38_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n27), .I3(GND_net), .O(n5571));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_75 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [12]), .I3(fifo_data_out[12]), .O(n10578));
    defparam i12_4_lut_4_lut_adj_75.LUT_INIT = 16'h3120;
    SB_LUT4 i4283_3_lut (.I0(\REG.mem_44_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n21), .I3(GND_net), .O(n5666));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4635_3_lut (.I0(\REG.mem_63_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n2), .I3(GND_net), .O(n6018));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4189_3_lut (.I0(\REG.mem_38_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n27), .I3(GND_net), .O(n5572));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4285_3_lut (.I0(\REG.mem_44_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n21), .I3(GND_net), .O(n5668));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4190_3_lut (.I0(\REG.mem_39_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n26), .I3(GND_net), .O(n5573));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4286_3_lut (.I0(\REG.mem_44_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n21), .I3(GND_net), .O(n5669));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4702_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [0]), .I3(fifo_data_out[0]), .O(n6085));
    defparam i4702_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4287_3_lut (.I0(\REG.mem_44_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n21), .I3(GND_net), .O(n5670));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4636_3_lut (.I0(\REG.mem_63_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n2), .I3(GND_net), .O(n6019));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4213_3_lut (.I0(\REG.mem_40_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n25), .I3(GND_net), .O(n5596));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4192_3_lut (.I0(\REG.mem_39_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n26), .I3(GND_net), .O(n5575));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4193_3_lut (.I0(\REG.mem_39_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n26), .I3(GND_net), .O(n5576));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_76 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [11]), .I3(fifo_data_out[11]), .O(n10576));
    defparam i12_4_lut_4_lut_adj_76.LUT_INIT = 16'h3120;
    SB_LUT4 i4194_3_lut (.I0(\REG.mem_39_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n26), .I3(GND_net), .O(n5577));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3516_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4899));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i3516_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4195_3_lut (.I0(\REG.mem_39_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n26), .I3(GND_net), .O(n5578));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4196_3_lut (.I0(\REG.mem_39_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n26), .I3(GND_net), .O(n5579));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4197_3_lut (.I0(\REG.mem_39_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n26), .I3(GND_net), .O(n5580));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3514_3_lut (.I0(rx_buf_byte[0]), .I1(rx_shift_reg[0]), .I2(n3495), 
            .I3(GND_net), .O(n4897));   // src/spi.v(76[8] 221[4])
    defparam i3514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4288_3_lut (.I0(\REG.mem_44_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n21), .I3(GND_net), .O(n5671));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_77 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [10]), .I3(fifo_data_out[10]), .O(n10574));
    defparam i12_4_lut_4_lut_adj_77.LUT_INIT = 16'h3120;
    SB_LUT4 i4738_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [2]), .I3(fifo_data_out[2]), .O(n6121));
    defparam i4738_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4637_3_lut (.I0(\REG.mem_63_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n2), .I3(GND_net), .O(n6020));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4290_3_lut (.I0(\REG.mem_45_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n20), .I3(GND_net), .O(n5673));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4291_3_lut (.I0(\REG.mem_45_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n20), .I3(GND_net), .O(n5674));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4292_3_lut (.I0(\REG.mem_45_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n20), .I3(GND_net), .O(n5675));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3539_4_lut (.I0(RESET_c), .I1(rd_addr_r_adj_121[2]), .I2(rd_addr_p1_w_adj_123[2]), 
            .I3(empty_o_N_1149), .O(n4922));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i3539_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i4109_3_lut (.I0(\REG.mem_35_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n30), .I3(GND_net), .O(n5492));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4293_3_lut (.I0(\REG.mem_45_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n20), .I3(GND_net), .O(n5676));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3520_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4903));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i3520_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4110_3_lut (.I0(\REG.mem_35_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n30), .I3(GND_net), .O(n5493));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4294_3_lut (.I0(\REG.mem_45_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n20), .I3(GND_net), .O(n5677));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3521_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4904));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i3521_2_lut.LUT_INIT = 16'h4444;
    SB_DFF tx_data_byte_r_i0_i7 (.Q(tx_data_byte[7]), .C(SLM_CLK_c), .D(n4942));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 i3524_2_lut (.I0(n2352), .I1(DEBUG_8_c_0_c), .I2(GND_net), 
            .I3(GND_net), .O(n4907));   // src/usb3_if.v(88[8] 191[4])
    defparam i3524_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3526_2_lut (.I0(uart_rx_complete_prev), .I1(debug_led3), .I2(GND_net), 
            .I3(GND_net), .O(n4909));   // src/top.v(1065[8] 1071[4])
    defparam i3526_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3527_2_lut (.I0(reset_per_frame_latched), .I1(n571), .I2(GND_net), 
            .I3(GND_net), .O(n4910));   // src/usb3_if.v(98[9] 189[16])
    defparam i3527_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4295_3_lut (.I0(\REG.mem_45_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n20), .I3(GND_net), .O(n5678));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4214_3_lut (.I0(\REG.mem_40_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n25), .I3(GND_net), .O(n5597));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4638_3_lut (.I0(\REG.mem_63_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n2), .I3(GND_net), .O(n6021));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4111_3_lut (.I0(\REG.mem_35_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n30), .I3(GND_net), .O(n5494));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4215_3_lut (.I0(\REG.mem_40_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n25), .I3(GND_net), .O(n5598));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4215_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF fifo_write_cmd_79 (.Q(fifo_write_cmd), .C(SLM_CLK_c), .D(n4939));   // src/top.v(889[8] 898[4])
    SB_LUT4 i4216_3_lut (.I0(\REG.mem_40_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n25), .I3(GND_net), .O(n5599));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_78 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [15]), .I3(fifo_data_out[15]), .O(n10588));
    defparam i12_4_lut_4_lut_adj_78.LUT_INIT = 16'h3120;
    SB_LUT4 i4112_3_lut (.I0(\REG.mem_35_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n30), .I3(GND_net), .O(n5495));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4217_3_lut (.I0(\REG.mem_40_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n25), .I3(GND_net), .O(n5600));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4113_3_lut (.I0(\REG.mem_35_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n30), .I3(GND_net), .O(n5496));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4296_3_lut (.I0(\REG.mem_45_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n20), .I3(GND_net), .O(n5679));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4297_3_lut (.I0(\REG.mem_45_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n20), .I3(GND_net), .O(n5680));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4114_3_lut (.I0(\REG.mem_35_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n30), .I3(GND_net), .O(n5497));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4218_3_lut (.I0(\REG.mem_40_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n25), .I3(GND_net), .O(n5601));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4115_3_lut (.I0(\REG.mem_35_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n30), .I3(GND_net), .O(n5498));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4298_3_lut (.I0(\REG.mem_45_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n20), .I3(GND_net), .O(n5681));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4219_3_lut (.I0(\REG.mem_40_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n25), .I3(GND_net), .O(n5602));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4219_3_lut.LUT_INIT = 16'hcaca;
=======
    SB_LUT4 i4787_3_lut (.I0(\REG.mem_20_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n13), .I3(GND_net), .O(n6261));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4788_3_lut (.I0(\REG.mem_20_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n13), .I3(GND_net), .O(n6262));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5487_3_lut (.I0(r_Tx_Data[2]), .I1(fifo_temp_output[2]), .I2(n4314), 
            .I3(GND_net), .O(n6961));   // src/uart_tx.v(38[10] 141[8])
    defparam i5487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4977_3_lut (.I0(\REG.mem_26_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n7), .I3(GND_net), .O(n6451));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4978_3_lut (.I0(\REG.mem_26_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n7), .I3(GND_net), .O(n6452));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4789_3_lut (.I0(\REG.mem_20_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n13), .I3(GND_net), .O(n6263));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5488_3_lut (.I0(r_Tx_Data[3]), .I1(fifo_temp_output[3]), .I2(n4314), 
            .I3(GND_net), .O(n6962));   // src/uart_tx.v(38[10] 141[8])
    defparam i5488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4979_3_lut (.I0(\REG.mem_26_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n7), .I3(GND_net), .O(n6453));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4790_3_lut (.I0(\REG.mem_20_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n13), .I3(GND_net), .O(n6264));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4980_3_lut (.I0(\REG.mem_26_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n7), .I3(GND_net), .O(n6454));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5489_3_lut (.I0(r_Tx_Data[4]), .I1(fifo_temp_output[4]), .I2(n4314), 
            .I3(GND_net), .O(n6963));   // src/uart_tx.v(38[10] 141[8])
    defparam i5489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4791_3_lut (.I0(\REG.mem_20_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n13), .I3(GND_net), .O(n6265));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4792_3_lut (.I0(\REG.mem_20_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n13), .I3(GND_net), .O(n6266));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4981_3_lut (.I0(\REG.mem_26_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n7), .I3(GND_net), .O(n6455));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4982_3_lut (.I0(\REG.mem_26_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n7), .I3(GND_net), .O(n6456));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4793_3_lut (.I0(\REG.mem_20_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n13), .I3(GND_net), .O(n6267));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5490_3_lut (.I0(r_Tx_Data[5]), .I1(fifo_temp_output[5]), .I2(n4314), 
            .I3(GND_net), .O(n6964));   // src/uart_tx.v(38[10] 141[8])
    defparam i5490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4794_3_lut (.I0(\REG.mem_20_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n13), .I3(GND_net), .O(n6268));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4983_3_lut (.I0(\REG.mem_26_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n7), .I3(GND_net), .O(n6457));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10870_2_lut (.I0(tx_data_byte[2]), .I1(tx_data_byte[4]), .I2(GND_net), 
            .I3(GND_net), .O(n12978));
    defparam i10870_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10941_4_lut (.I0(tx_data_byte[3]), .I1(tx_data_byte[7]), .I2(tx_data_byte[5]), 
            .I3(n12978), .O(n13052));
    defparam i10941_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i12303_4_lut (.I0(tx_data_byte[0]), .I1(tx_data_byte[1]), .I2(tx_data_byte[6]), 
            .I3(n13052), .O(multi_byte_spi_trans_flag_r_N_72));   // src/top.v(1214[10:31])
    defparam i12303_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i4984_3_lut (.I0(\REG.mem_26_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n7), .I3(GND_net), .O(n6458));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5491_3_lut (.I0(r_Tx_Data[6]), .I1(fifo_temp_output[6]), .I2(n4314), 
            .I3(GND_net), .O(n6965));   // src/uart_tx.v(38[10] 141[8])
    defparam i5491_3_lut.LUT_INIT = 16'hcaca;
>>>>>>> Stashed changes
>>>>>>> master
    SB_IO CTS_pad (.PACKAGE_PIN(CTS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CTS_pad.PIN_TYPE = 6'b011001;
    defparam CTS_pad.PULLUP = 1'b0;
    defparam CTS_pad.NEG_TRIGGER = 1'b0;
    defparam CTS_pad.IO_STANDARD = "SB_LVCMOS";
<<<<<<< HEAD
    SB_LUT4 i4173_2_lut (.I0(is_tx_fifo_full_flag), .I1(spi_rx_byte_ready), 
            .I2(GND_net), .I3(GND_net), .O(n5632));   // src/top.v(980[8] 989[4])
    defparam i4173_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4175_4_lut (.I0(\REG.mem_3_0 ), .I1(DEBUG_3_c_0), .I2(n27), 
            .I3(wr_addr_r[4]), .O(n5634));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4175_4_lut.LUT_INIT = 16'haaca;
    SB_DFF tx_data_byte_r_i0_i2 (.Q(tx_data_byte[2]), .C(SLM_CLK_c), .D(n5724));   // src/top.v(1165[8] 1232[4])
    SB_LUT4 i4176_4_lut (.I0(\REG.mem_4_0 ), .I1(DEBUG_3_c_0), .I2(n29), 
            .I3(wr_addr_r[4]), .O(n5635));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4176_4_lut.LUT_INIT = 16'haaca;
    SB_DFF reset_all_r_77 (.Q(reset_all_w), .C(SLM_CLK_c), .D(reset_all_w_N_61));   // src/top.v(246[8] 264[4])
    SB_LUT4 i4250_4_lut (.I0(pc_data_rx[7]), .I1(r_Rx_Data), .I2(n6690), 
            .I3(n8012), .O(n5709));   // src/uart_rx.v(49[10] 144[8])
    defparam i4250_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i4251_3_lut (.I0(r_Tx_Data[7]), .I1(fifo_temp_output[7]), .I2(n4715), 
            .I3(GND_net), .O(n5710));   // src/uart_tx.v(38[10] 141[8])
    defparam i4251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4252_3_lut (.I0(r_Tx_Data[6]), .I1(fifo_temp_output[6]), .I2(n4715), 
            .I3(GND_net), .O(n5711));   // src/uart_tx.v(38[10] 141[8])
    defparam i4252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4253_3_lut (.I0(r_Tx_Data[5]), .I1(fifo_temp_output[5]), .I2(n4715), 
            .I3(GND_net), .O(n5712));   // src/uart_tx.v(38[10] 141[8])
    defparam i4253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4178_4_lut (.I0(\REG.mem_5_0 ), .I1(DEBUG_3_c_0), .I2(n31), 
            .I3(wr_addr_r[4]), .O(n5637));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4178_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i4179_4_lut (.I0(\REG.mem_6_0 ), .I1(DEBUG_3_c_0), .I2(n33), 
            .I3(wr_addr_r[4]), .O(n5638));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4179_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 led_counter_1344_1403_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(DEBUG_0_c_24), .I3(n10373), .O(n106_adj_1406)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4180_4_lut (.I0(\REG.mem_7_0 ), .I1(DEBUG_3_c_0), .I2(n35), 
            .I3(wr_addr_r[4]), .O(n5639));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4180_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i4254_3_lut (.I0(r_Tx_Data[4]), .I1(fifo_temp_output[4]), .I2(n4715), 
            .I3(GND_net), .O(n5713));   // src/uart_tx.v(38[10] 141[8])
    defparam i4254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1344_1403_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n2), .I3(n10372), .O(n107)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1344_1403_add_4_25 (.CI(n10372), .I0(GND_net), 
            .I1(n2), .CO(n10373));
    SB_LUT4 led_counter_1344_1403_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_1411), .I3(n10371), .O(n108)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1344_1403_add_4_24 (.CI(n10371), .I0(GND_net), 
            .I1(n3_adj_1411), .CO(n10372));
    SB_LUT4 led_counter_1344_1403_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_1418), .I3(n10370), .O(n109)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4255_3_lut (.I0(r_Tx_Data[3]), .I1(fifo_temp_output[3]), .I2(n4715), 
            .I3(GND_net), .O(n5714));   // src/uart_tx.v(38[10] 141[8])
    defparam i4255_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1344_1403_add_4_23 (.CI(n10370), .I0(GND_net), 
            .I1(n4_adj_1418), .CO(n10371));
    SB_LUT4 led_counter_1344_1403_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5), .I3(n10369), .O(n110)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_22_lut.LUT_INIT = 16'hC33C;
=======
<<<<<<< Updated upstream
    SB_CARRY led_counter_1186_1260_add_4_6 (.CI(n10175), .I0(GND_net), .I1(n21_adj_66), 
            .CO(n10176));
    SB_LUT4 i4299_3_lut (.I0(\REG.mem_45_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n20), .I3(GND_net), .O(n5682));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4299_3_lut.LUT_INIT = 16'hcaca;
=======
    SB_LUT4 i4985_3_lut (.I0(\REG.mem_26_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n7), .I3(GND_net), .O(n6459));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4986_3_lut (.I0(\REG.mem_26_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n7), .I3(GND_net), .O(n6460));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4795_3_lut (.I0(\REG.mem_20_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n13), .I3(GND_net), .O(n6269));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4987_3_lut (.I0(\REG.mem_26_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n7), .I3(GND_net), .O(n6461));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4796_3_lut (.I0(\REG.mem_21_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n12), .I3(GND_net), .O(n6270));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4797_3_lut (.I0(\REG.mem_21_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n12), .I3(GND_net), .O(n6271));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4988_3_lut (.I0(\REG.mem_27_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n6), .I3(GND_net), .O(n6462));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5492_3_lut (.I0(r_Tx_Data[7]), .I1(fifo_temp_output[7]), .I2(n4314), 
            .I3(GND_net), .O(n6966));   // src/uart_tx.v(38[10] 141[8])
    defparam i5492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4989_3_lut (.I0(\REG.mem_27_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n6), .I3(GND_net), .O(n6463));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4990_3_lut (.I0(\REG.mem_27_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n6), .I3(GND_net), .O(n6464));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4991_3_lut (.I0(\REG.mem_27_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n6), .I3(GND_net), .O(n6465));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4992_3_lut (.I0(\REG.mem_27_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n6), .I3(GND_net), .O(n6466));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4993_3_lut (.I0(\REG.mem_27_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n6), .I3(GND_net), .O(n6467));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4994_3_lut (.I0(\REG.mem_27_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n6), .I3(GND_net), .O(n6468));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4798_3_lut (.I0(\REG.mem_21_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n12), .I3(GND_net), .O(n6272));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4995_3_lut (.I0(\REG.mem_27_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n6), .I3(GND_net), .O(n6469));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 reset_all_w_I_0_1_lut (.I0(reset_all_w), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(RESET_c));   // src/top.v(295[16:28])
    defparam reset_all_w_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4799_3_lut (.I0(\REG.mem_21_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n12), .I3(GND_net), .O(n6273));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4800_3_lut (.I0(\REG.mem_21_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n12), .I3(GND_net), .O(n6274));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4996_3_lut (.I0(\REG.mem_27_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n6), .I3(GND_net), .O(n6470));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4997_3_lut (.I0(\REG.mem_27_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n6), .I3(GND_net), .O(n6471));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5493_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[0]), .I2(n4_adj_1435), 
            .I3(n4790), .O(n6967));   // src/uart_rx.v(49[10] 144[8])
    defparam i5493_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4998_3_lut (.I0(\REG.mem_27_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n6), .I3(GND_net), .O(n6472));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4999_3_lut (.I0(\REG.mem_27_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n6), .I3(GND_net), .O(n6473));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut (.I0(tx_shift_reg[0]), .I1(n2407), .I2(n4837), .I3(tx_data_byte[0]), 
            .O(n12537));   // src/spi.v(76[8] 221[4])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i5000_3_lut (.I0(\REG.mem_27_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n6), .I3(GND_net), .O(n6474));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5001_3_lut (.I0(\REG.mem_27_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n6), .I3(GND_net), .O(n6475));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4801_3_lut (.I0(\REG.mem_21_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n12), .I3(GND_net), .O(n6275));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4802_3_lut (.I0(\REG.mem_21_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n12), .I3(GND_net), .O(n6276));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5002_3_lut (.I0(\REG.mem_27_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n6), .I3(GND_net), .O(n6476));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5003_3_lut (.I0(\REG.mem_27_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n6), .I3(GND_net), .O(n6477));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10831_4_lut (.I0(n4446), .I1(fifo_read_cmd), .I2(wr_addr_r_adj_1517[1]), 
            .I3(rd_addr_r_adj_1520[1]), .O(n12938));
    defparam i10831_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i5004_3_lut (.I0(\REG.mem_27_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n6), .I3(GND_net), .O(n6478));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4803_3_lut (.I0(\REG.mem_21_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n12), .I3(GND_net), .O(n6277));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4804_3_lut (.I0(\REG.mem_21_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n12), .I3(GND_net), .O(n6278));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4805_3_lut (.I0(\REG.mem_21_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n12), .I3(GND_net), .O(n6279));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5005_3_lut (.I0(\REG.mem_27_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n6), .I3(GND_net), .O(n6479));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4806_3_lut (.I0(\REG.mem_21_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n12), .I3(GND_net), .O(n6280));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5006_3_lut (.I0(\REG.mem_27_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n6), .I3(GND_net), .O(n6480));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(reset_all_w), .I1(n15), .I2(wr_fifo_en_w_adj_1416), 
            .I3(n12215), .O(n12439));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut.LUT_INIT = 16'h5444;
    SB_LUT4 i5007_3_lut (.I0(\REG.mem_27_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n6), .I3(GND_net), .O(n6481));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5501_3_lut (.I0(rx_shift_reg[1]), .I1(rx_shift_reg[0]), .I2(n4884), 
            .I3(GND_net), .O(n6975));   // src/spi.v(76[8] 221[4])
    defparam i5501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4807_3_lut (.I0(\REG.mem_21_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n12), .I3(GND_net), .O(n6281));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5008_3_lut (.I0(\REG.mem_27_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n6), .I3(GND_net), .O(n6482));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5502_3_lut (.I0(rx_shift_reg[2]), .I1(rx_shift_reg[1]), .I2(n4884), 
            .I3(GND_net), .O(n6976));   // src/spi.v(76[8] 221[4])
    defparam i5502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5009_3_lut (.I0(\REG.mem_27_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n6), .I3(GND_net), .O(n6483));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5010_3_lut (.I0(\REG.mem_27_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n6), .I3(GND_net), .O(n6484));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5011_3_lut (.I0(\REG.mem_27_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n6), .I3(GND_net), .O(n6485));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4808_3_lut (.I0(\REG.mem_21_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n12), .I3(GND_net), .O(n6282));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5012_3_lut (.I0(\REG.mem_27_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n6), .I3(GND_net), .O(n6486));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5503_3_lut (.I0(rx_shift_reg[3]), .I1(rx_shift_reg[2]), .I2(n4884), 
            .I3(GND_net), .O(n6977));   // src/spi.v(76[8] 221[4])
    defparam i5503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4809_3_lut (.I0(\REG.mem_21_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n12), .I3(GND_net), .O(n6283));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5013_3_lut (.I0(\REG.mem_27_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n6), .I3(GND_net), .O(n6487));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5014_3_lut (.I0(\REG.mem_27_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n6), .I3(GND_net), .O(n6488));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5504_3_lut (.I0(rx_shift_reg[4]), .I1(rx_shift_reg[3]), .I2(n4884), 
            .I3(GND_net), .O(n6978));   // src/spi.v(76[8] 221[4])
    defparam i5504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5505_3_lut (.I0(rx_shift_reg[5]), .I1(rx_shift_reg[4]), .I2(n4884), 
            .I3(GND_net), .O(n6979));   // src/spi.v(76[8] 221[4])
    defparam i5505_3_lut.LUT_INIT = 16'hcaca;
>>>>>>> Stashed changes
>>>>>>> master
    SB_IO DTR_pad (.PACKAGE_PIN(DTR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DTR_pad.PIN_TYPE = 6'b011001;
    defparam DTR_pad.PULLUP = 1'b0;
    defparam DTR_pad.NEG_TRIGGER = 1'b0;
    defparam DTR_pad.IO_STANDARD = "SB_LVCMOS";
<<<<<<< HEAD
    SB_LUT4 i4366_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[0]), .I2(n4_adj_1413), 
            .I3(n5019), .O(n5825));   // src/uart_rx.v(49[10] 144[8])
    defparam i4366_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY led_counter_1344_1403_add_4_22 (.CI(n10369), .I0(GND_net), 
            .I1(n5), .CO(n10370));
    SB_LUT4 led_counter_1344_1403_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_1408), .I3(n10368), .O(n111)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_21_lut.LUT_INIT = 16'hC33C;
=======
<<<<<<< Updated upstream
    SB_LUT4 i4116_3_lut (.I0(\REG.mem_35_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n30), .I3(GND_net), .O(n5499));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4116_3_lut.LUT_INIT = 16'hcaca;
=======
    SB_LUT4 i5015_3_lut (.I0(\REG.mem_27_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n6), .I3(GND_net), .O(n6489));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4810_3_lut (.I0(\REG.mem_21_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n12), .I3(GND_net), .O(n6284));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4811_3_lut (.I0(\REG.mem_21_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n12), .I3(GND_net), .O(n6285));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5016_3_lut (.I0(\REG.mem_27_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n6), .I3(GND_net), .O(n6490));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5017_3_lut (.I0(\REG.mem_27_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n6), .I3(GND_net), .O(n6491));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5506_3_lut (.I0(rx_shift_reg[6]), .I1(rx_shift_reg[5]), .I2(n4884), 
            .I3(GND_net), .O(n6980));   // src/spi.v(76[8] 221[4])
    defparam i5506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5018_3_lut (.I0(\REG.mem_27_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n6), .I3(GND_net), .O(n6492));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4812_3_lut (.I0(\REG.mem_21_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n12), .I3(GND_net), .O(n6286));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5507_3_lut (.I0(rx_shift_reg[7]), .I1(rx_shift_reg[6]), .I2(n4884), 
            .I3(GND_net), .O(n6981));   // src/spi.v(76[8] 221[4])
    defparam i5507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4813_3_lut (.I0(\REG.mem_21_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n12), .I3(GND_net), .O(n6287));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4814_3_lut (.I0(\REG.mem_21_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n12), .I3(GND_net), .O(n6288));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5508_3_lut (.I0(rx_buf_byte[1]), .I1(rx_shift_reg[1]), .I2(n3963), 
            .I3(GND_net), .O(n6982));   // src/spi.v(76[8] 221[4])
    defparam i5508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4815_3_lut (.I0(\REG.mem_21_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n12), .I3(GND_net), .O(n6289));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5019_3_lut (.I0(\REG.mem_27_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n6), .I3(GND_net), .O(n6493));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4816_3_lut (.I0(\REG.mem_21_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n12), .I3(GND_net), .O(n6290));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5509_3_lut (.I0(rx_buf_byte[2]), .I1(rx_shift_reg[2]), .I2(n3963), 
            .I3(GND_net), .O(n6983));   // src/spi.v(76[8] 221[4])
    defparam i5509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4817_3_lut (.I0(\REG.mem_21_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n12), .I3(GND_net), .O(n6291));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4818_3_lut (.I0(\REG.mem_21_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n12), .I3(GND_net), .O(n6292));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4819_3_lut (.I0(\REG.mem_21_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n12), .I3(GND_net), .O(n6293));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4820_3_lut (.I0(\REG.mem_21_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n12), .I3(GND_net), .O(n6294));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4821_3_lut (.I0(\REG.mem_21_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n12), .I3(GND_net), .O(n6295));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4822_3_lut (.I0(\REG.mem_21_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n12), .I3(GND_net), .O(n6296));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5510_3_lut (.I0(rx_buf_byte[3]), .I1(rx_shift_reg[3]), .I2(n3963), 
            .I3(GND_net), .O(n6984));   // src/spi.v(76[8] 221[4])
    defparam i5510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4823_3_lut (.I0(\REG.mem_21_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n12), .I3(GND_net), .O(n6297));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4823_3_lut.LUT_INIT = 16'hcaca;
>>>>>>> Stashed changes
>>>>>>> master
    SB_IO DSR_pad (.PACKAGE_PIN(DSR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DSR_pad.PIN_TYPE = 6'b011001;
    defparam DSR_pad.PULLUP = 1'b0;
    defparam DSR_pad.NEG_TRIGGER = 1'b0;
    defparam DSR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DCD_pad (.PACKAGE_PIN(DCD), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DCD_pad.PIN_TYPE = 6'b011001;
    defparam DCD_pad.PULLUP = 1'b0;
    defparam DCD_pad.NEG_TRIGGER = 1'b0;
    defparam DCD_pad.IO_STANDARD = "SB_LVCMOS";
<<<<<<< HEAD
    SB_IO UART_TX_pad (.PACKAGE_PIN(UART_TX), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(UART_TX_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UART_TX_pad.PIN_TYPE = 6'b011001;
    defparam UART_TX_pad.PULLUP = 1'b0;
    defparam UART_TX_pad.NEG_TRIGGER = 1'b0;
    defparam UART_TX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY led_counter_1344_1403_add_4_21 (.CI(n10368), .I0(GND_net), 
            .I1(n6_adj_1408), .CO(n10369));
    SB_LUT4 i1982_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n3426));   // src/top.v(1165[8] 1232[4])
    defparam i1982_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 led_counter_1344_1403_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_1412), .I3(n10367), .O(n112)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_DFF tx_data_byte_r_i0_i3 (.Q(tx_data_byte[3]), .C(SLM_CLK_c), .D(n5720));   // src/top.v(1165[8] 1232[4])
    SB_CARRY led_counter_1344_1403_add_4_20 (.CI(n10367), .I0(GND_net), 
            .I1(n7_adj_1412), .CO(n10368));
    SB_LUT4 led_counter_1344_1403_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8), .I3(n10366), .O(n113)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1344_1403_add_4_19 (.CI(n10366), .I0(GND_net), 
            .I1(n8), .CO(n10367));
    SB_LUT4 led_counter_1344_1403_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9), .I3(n10365), .O(n114)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1344_1403_add_4_18 (.CI(n10365), .I0(GND_net), 
            .I1(n9), .CO(n10366));
    SB_LUT4 led_counter_1344_1403_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10), .I3(n10364), .O(n115)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n5101), 
            .I3(debug_led3), .O(n10608));   // src/uart_rx.v(49[10] 144[8])
=======
<<<<<<< Updated upstream
    SB_LUT4 i4118_3_lut (.I0(\REG.mem_35_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n30), .I3(GND_net), .O(n5501));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4118_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DEBUG_8_c_0_pad (.PACKAGE_PIN(FIFO_D0), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(DEBUG_8_c_0_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_8_c_0_pad.PIN_TYPE = 6'b000001;
    defparam DEBUG_8_c_0_pad.PULLUP = 1'b0;
    defparam DEBUG_8_c_0_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_8_c_0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4220_3_lut (.I0(\REG.mem_40_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n25), .I3(GND_net), .O(n5603));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4221_3_lut (.I0(\REG.mem_40_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n25), .I3(GND_net), .O(n5604));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_79 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [4]), .I3(fifo_data_out[4]), .O(n10562));
    defparam i12_4_lut_4_lut_adj_79.LUT_INIT = 16'h3120;
    SB_LUT4 i4300_3_lut (.I0(\REG.mem_45_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n20), .I3(GND_net), .O(n5683));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4301_3_lut (.I0(\REG.mem_45_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n20), .I3(GND_net), .O(n5684));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4119_3_lut (.I0(\REG.mem_35_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n30), .I3(GND_net), .O(n5502));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4302_3_lut (.I0(\REG.mem_45_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n20), .I3(GND_net), .O(n5685));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4641_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[5]), .I2(GND_net), 
            .I3(GND_net), .O(n6024));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4641_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4303_3_lut (.I0(\REG.mem_45_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n20), .I3(GND_net), .O(n5686));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4222_3_lut (.I0(\REG.mem_40_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n25), .I3(GND_net), .O(n5605));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4223_3_lut (.I0(\REG.mem_41_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5606));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_80 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [8]), .I3(fifo_data_out[8]), .O(n10570));
    defparam i12_4_lut_4_lut_adj_80.LUT_INIT = 16'h3120;
    SB_LUT4 i4304_3_lut (.I0(\REG.mem_45_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n20), .I3(GND_net), .O(n5687));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4224_3_lut (.I0(\REG.mem_41_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5607));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4225_3_lut (.I0(\REG.mem_41_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5608));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_81 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [6]), .I3(fifo_data_out[6]), .O(n10566));
    defparam i12_4_lut_4_lut_adj_81.LUT_INIT = 16'h3120;
    SB_LUT4 i4120_3_lut (.I0(\REG.mem_35_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n30), .I3(GND_net), .O(n5503));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4305_3_lut (.I0(\REG.mem_45_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n20), .I3(GND_net), .O(n5688));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4735_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [1]), .I3(fifo_data_out[1]), .O(n6118));
    defparam i4735_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4306_3_lut (.I0(\REG.mem_46_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n19), .I3(GND_net), .O(n5689));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4226_3_lut (.I0(\REG.mem_41_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5609));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4307_3_lut (.I0(\REG.mem_46_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n19), .I3(GND_net), .O(n5690));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_82 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [7]), .I3(fifo_data_out[7]), .O(n10568));
    defparam i12_4_lut_4_lut_adj_82.LUT_INIT = 16'h3120;
    SB_LUT4 i4227_3_lut (.I0(\REG.mem_41_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5610));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4228_3_lut (.I0(\REG.mem_41_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5611));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4308_3_lut (.I0(\REG.mem_46_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n19), .I3(GND_net), .O(n5691));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4309_3_lut (.I0(\REG.mem_46_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n19), .I3(GND_net), .O(n5692));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4121_3_lut (.I0(\REG.mem_35_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n30), .I3(GND_net), .O(n5504));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4122_3_lut (.I0(\REG.mem_35_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n30), .I3(GND_net), .O(n5505));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4310_3_lut (.I0(\REG.mem_46_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n19), .I3(GND_net), .O(n5693));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3528_2_lut (.I0(reset_per_frame_latched), .I1(n575), .I2(GND_net), 
            .I3(GND_net), .O(n4911));   // src/usb3_if.v(98[9] 189[16])
    defparam i3528_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4123_3_lut (.I0(\REG.mem_35_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n30), .I3(GND_net), .O(n5506));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4229_3_lut (.I0(\REG.mem_41_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5612));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4311_3_lut (.I0(\REG.mem_46_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n19), .I3(GND_net), .O(n5694));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4312_3_lut (.I0(\REG.mem_46_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n19), .I3(GND_net), .O(n5695));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4313_3_lut (.I0(\REG.mem_46_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n19), .I3(GND_net), .O(n5696));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4314_3_lut (.I0(\REG.mem_46_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n19), .I3(GND_net), .O(n5697));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4314_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i0 (.Q(n25_adj_62), .C(SLM_CLK_c), .D(n130));   // src/top.v(203[20:35])
    SB_LUT4 i4315_3_lut (.I0(\REG.mem_46_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n19), .I3(GND_net), .O(n5698));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_83 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [3]), .I3(fifo_data_out[3]), .O(n10556));
    defparam i12_4_lut_4_lut_adj_83.LUT_INIT = 16'h3120;
    SB_LUT4 i4316_3_lut (.I0(\REG.mem_46_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n19), .I3(GND_net), .O(n5699));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_84 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [5]), .I3(fifo_data_out[5]), .O(n10564));
    defparam i12_4_lut_4_lut_adj_84.LUT_INIT = 16'h3120;
    SB_LUT4 i4124_3_lut (.I0(\REG.mem_35_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n30), .I3(GND_net), .O(n5507));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4317_3_lut (.I0(\REG.mem_46_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n19), .I3(GND_net), .O(n5700));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4318_3_lut (.I0(\REG.mem_46_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n19), .I3(GND_net), .O(n5701));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4318_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_clk_counter_i3_1187__i3 (.Q(reset_clk_counter[3]), .C(SLM_CLK_c), 
           .D(n10293));   // src/top.v(259[27:51])
    SB_LUT4 i12_4_lut_4_lut_adj_85 (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [9]), .I3(fifo_data_out[9]), .O(n10572));
    defparam i12_4_lut_4_lut_adj_85.LUT_INIT = 16'h3120;
    SB_LUT4 i4230_3_lut (.I0(\REG.mem_41_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5613));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4319_3_lut (.I0(\REG.mem_46_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n19), .I3(GND_net), .O(n5702));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4231_3_lut (.I0(\REG.mem_41_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5614));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4232_3_lut (.I0(\REG.mem_41_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5615));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3540_3_lut (.I0(tx_addr_byte[0]), .I1(tx_data_byte[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4923));   // src/top.v(1074[8] 1141[4])
    defparam i3540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4233_3_lut (.I0(\REG.mem_41_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5616));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4234_3_lut (.I0(\REG.mem_41_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5617));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4320_3_lut (.I0(\REG.mem_46_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n19), .I3(GND_net), .O(n5703));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4235_3_lut (.I0(\REG.mem_41_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5618));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4321_3_lut (.I0(\REG.mem_46_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n19), .I3(GND_net), .O(n5704));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4321_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_clk_counter_i3_1187__i2 (.Q(reset_clk_counter[2]), .C(SLM_CLK_c), 
           .D(n10295));   // src/top.v(259[27:51])
    SB_DFF reset_clk_counter_i3_1187__i1 (.Q(reset_clk_counter[1]), .C(SLM_CLK_c), 
           .D(n10291));   // src/top.v(259[27:51])
    SB_DFF led_counter_1186_1260__i24 (.Q(DEBUG_0_c_24), .C(SLM_CLK_c), 
           .D(n106));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i23 (.Q(n2_adj_75), .C(SLM_CLK_c), .D(n107));   // src/top.v(203[20:35])
    SB_LUT4 i4236_3_lut (.I0(\REG.mem_41_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5619));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4236_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i22 (.Q(n3), .C(SLM_CLK_c), .D(n108));   // src/top.v(203[20:35])
    SB_LUT4 i4237_3_lut (.I0(\REG.mem_41_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5620));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4237_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i21 (.Q(n4_adj_74), .C(SLM_CLK_c), .D(n109));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i20 (.Q(n5), .C(SLM_CLK_c), .D(n110));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i19 (.Q(n6), .C(SLM_CLK_c), .D(n111));   // src/top.v(203[20:35])
    SB_LUT4 i4322_3_lut (.I0(\REG.mem_47_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n18), .I3(GND_net), .O(n5705));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4323_3_lut (.I0(\REG.mem_47_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n18), .I3(GND_net), .O(n5706));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4324_3_lut (.I0(\REG.mem_47_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n18), .I3(GND_net), .O(n5707));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4238_3_lut (.I0(\REG.mem_41_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n24_adj_61), .I3(GND_net), .O(n5621));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4325_3_lut (.I0(\REG.mem_47_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n18), .I3(GND_net), .O(n5708));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4239_3_lut (.I0(\REG.mem_42_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n23), .I3(GND_net), .O(n5622));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4326_3_lut (.I0(\REG.mem_47_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n18), .I3(GND_net), .O(n5709));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4326_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i18 (.Q(n7), .C(SLM_CLK_c), .D(n112));   // src/top.v(203[20:35])
    SB_LUT4 i4240_3_lut (.I0(\REG.mem_42_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n23), .I3(GND_net), .O(n5623));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4240_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i17 (.Q(n8_adj_73), .C(SLM_CLK_c), .D(n113));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i16 (.Q(n9), .C(SLM_CLK_c), .D(n114));   // src/top.v(203[20:35])
    SB_LUT4 i4241_3_lut (.I0(\REG.mem_42_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n23), .I3(GND_net), .O(n5624));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4241_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i15 (.Q(n10_adj_72), .C(SLM_CLK_c), .D(n115));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i14 (.Q(n11), .C(SLM_CLK_c), .D(n116));   // src/top.v(203[20:35])
    SB_LUT4 i4327_3_lut (.I0(\REG.mem_47_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n18), .I3(GND_net), .O(n5710));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4327_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i13 (.Q(n12), .C(SLM_CLK_c), .D(n117));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i12 (.Q(n13), .C(SLM_CLK_c), .D(n118));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i11 (.Q(n14), .C(SLM_CLK_c), .D(n119));   // src/top.v(203[20:35])
    SB_LUT4 i4242_3_lut (.I0(\REG.mem_42_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n23), .I3(GND_net), .O(n5625));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4242_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i10 (.Q(n15_adj_71), .C(SLM_CLK_c), .D(n120));   // src/top.v(203[20:35])
    SB_LUT4 i4243_3_lut (.I0(\REG.mem_42_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n23), .I3(GND_net), .O(n5626));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4243_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i9 (.Q(n16), .C(SLM_CLK_c), .D(n121));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i8 (.Q(n17_adj_70), .C(SLM_CLK_c), .D(n122));   // src/top.v(203[20:35])
    SB_LUT4 i4328_3_lut (.I0(\REG.mem_47_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n18), .I3(GND_net), .O(n5711));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4328_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i7 (.Q(n18_adj_69), .C(SLM_CLK_c), .D(n123));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i6 (.Q(n19_adj_68), .C(SLM_CLK_c), .D(n124));   // src/top.v(203[20:35])
    SB_LUT4 i4329_3_lut (.I0(\REG.mem_47_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n18), .I3(GND_net), .O(n5712));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4329_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i5 (.Q(n20_adj_67), .C(SLM_CLK_c), .D(n125));   // src/top.v(203[20:35])
    SB_LUT4 i4244_3_lut (.I0(\REG.mem_42_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n23), .I3(GND_net), .O(n5627));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4244_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i4 (.Q(n21_adj_66), .C(SLM_CLK_c), .D(n126));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i3 (.Q(n22_adj_65), .C(SLM_CLK_c), .D(n127));   // src/top.v(203[20:35])
    SB_LUT4 i4330_3_lut (.I0(\REG.mem_47_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n18), .I3(GND_net), .O(n5713));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4331_3_lut (.I0(\REG.mem_47_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n18), .I3(GND_net), .O(n5714));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_765[2]), 
            .I3(r_SM_Main[0]), .O(n4335));   // src/uart_rx.v(49[10] 144[8])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i4245_3_lut (.I0(\REG.mem_42_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n23), .I3(GND_net), .O(n5628));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4332_3_lut (.I0(\REG.mem_47_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n18), .I3(GND_net), .O(n5715));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4333_3_lut (.I0(\REG.mem_47_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n18), .I3(GND_net), .O(n5716));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4660_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[3]), .I2(GND_net), 
            .I3(GND_net), .O(n6043));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4660_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4334_3_lut (.I0(\REG.mem_47_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n18), .I3(GND_net), .O(n5717));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4334_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i2 (.Q(n23_adj_64), .C(SLM_CLK_c), .D(n128));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i1 (.Q(n24_adj_63), .C(SLM_CLK_c), .D(n129));   // src/top.v(203[20:35])
    SB_LUT4 i1_4_lut (.I0(rd_addr_r_adj_121[1]), .I1(rd_addr_r_adj_121[0]), 
            .I2(wr_addr_r_adj_118[1]), .I3(wr_addr_r_adj_118[0]), .O(n32));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut.LUT_INIT = 16'h8421;
    SB_LUT4 i4335_3_lut (.I0(\REG.mem_47_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n18), .I3(GND_net), .O(n5718));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4336_3_lut (.I0(\REG.mem_47_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n18), .I3(GND_net), .O(n5719));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n4335), 
            .I3(debug_led3), .O(n10406));   // src/uart_rx.v(49[10] 144[8])
>>>>>>> master
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_CARRY led_counter_1344_1403_add_4_17 (.CI(n10364), .I0(GND_net), 
            .I1(n10), .CO(n10365));
    SB_LUT4 i4256_3_lut (.I0(r_Tx_Data[2]), .I1(fifo_temp_output[2]), .I2(n4715), 
            .I3(GND_net), .O(n5715));   // src/uart_tx.v(38[10] 141[8])
    defparam i4256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1344_1403_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11), .I3(n10363), .O(n116)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1344_1403_add_4_16 (.CI(n10363), .I0(GND_net), 
            .I1(n11), .CO(n10364));
    SB_DFF even_byte_flag_89 (.Q(even_byte_flag), .C(SLM_CLK_c), .D(n3254));   // src/top.v(1165[8] 1232[4])
    SB_LUT4 led_counter_1344_1403_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12), .I3(n10362), .O(n117)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4257_3_lut (.I0(r_Tx_Data[1]), .I1(fifo_temp_output[1]), .I2(n4715), 
            .I3(GND_net), .O(n5716));   // src/uart_tx.v(38[10] 141[8])
    defparam i4257_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1344_1403_add_4_15 (.CI(n10362), .I0(GND_net), 
            .I1(n12), .CO(n10363));
    SB_LUT4 led_counter_1344_1403_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13), .I3(n10361), .O(n118)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1830_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n3254));   // src/top.v(1165[8] 1232[4])
    defparam i1830_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut (.I0(tx_shift_reg[0]), .I1(n2329), .I2(n5081), .I3(tx_data_byte[0]), 
            .O(n10792));   // src/spi.v(76[8] 221[4])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_IO FIFO_D0_pad (.PACKAGE_PIN(FIFO_D0), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D0_c_0));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D0_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D0_pad.PULLUP = 1'b0;
    defparam FIFO_D0_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY led_counter_1344_1403_add_4_14 (.CI(n10361), .I0(GND_net), 
            .I1(n13), .CO(n10362));
    SB_LUT4 led_counter_1344_1403_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14), .I3(n10360), .O(n119)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1344_1403_add_4_13 (.CI(n10360), .I0(GND_net), 
            .I1(n14), .CO(n10361));
    SB_LUT4 led_counter_1344_1403_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_1417), .I3(n10359), .O(n120)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1344_1403_add_4_12 (.CI(n10359), .I0(GND_net), 
            .I1(n15_adj_1417), .CO(n10360));
    SB_LUT4 led_counter_1344_1403_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16), .I3(n10358), .O(n121)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4181_4_lut (.I0(\REG.mem_8_0 ), .I1(DEBUG_3_c_0), .I2(n20), 
            .I3(wr_addr_r[4]), .O(n5640));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4181_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i4182_4_lut (.I0(\REG.mem_9_0 ), .I1(DEBUG_3_c_0), .I2(n22), 
            .I3(wr_addr_r[4]), .O(n5641));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4182_4_lut.LUT_INIT = 16'haaca;
    SB_CARRY led_counter_1344_1403_add_4_11 (.CI(n10358), .I0(GND_net), 
            .I1(n16), .CO(n10359));
    SB_LUT4 i4183_4_lut (.I0(\REG.mem_10_0 ), .I1(DEBUG_3_c_0), .I2(n24_adj_1404), 
            .I3(wr_addr_r[4]), .O(n5642));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4183_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i4258_4_lut (.I0(\REG.mem_21_0 ), .I1(DEBUG_3_c_0), .I2(n31), 
            .I3(wr_addr_r[4]), .O(n5717));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4258_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 led_counter_1344_1403_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17), .I3(n10357), .O(n122)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9662_4_lut (.I0(n1), .I1(fifo_read_cmd), .I2(wr_addr_r_adj_1490[1]), 
            .I3(rd_addr_r_adj_1493[1]), .O(n11239));
    defparam i9662_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i1_4_lut_adj_130 (.I0(RESET_c), .I1(n15), .I2(wr_fifo_en_w), 
            .I3(n10381), .O(n10640));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_adj_130.LUT_INIT = 16'ha888;
    SB_CARRY led_counter_1344_1403_add_4_10 (.CI(n10357), .I0(GND_net), 
            .I1(n17), .CO(n10358));
    SB_LUT4 led_counter_1344_1403_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18), .I3(n10356), .O(n123)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1344_1403_add_4_9 (.CI(n10356), .I0(GND_net), .I1(n18), 
            .CO(n10357));
    SB_LUT4 led_counter_1344_1403_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19), .I3(n10355), .O(n124)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1344_1403_add_4_8 (.CI(n10355), .I0(GND_net), .I1(n19), 
            .CO(n10356));
    SB_LUT4 led_counter_1344_1403_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_1416), .I3(n10354), .O(n125)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1344_1403_add_4_7 (.CI(n10354), .I0(GND_net), .I1(n20_adj_1416), 
            .CO(n10355));
    SB_LUT4 led_counter_1344_1403_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_1414), .I3(n10353), .O(n126)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1344_1403_add_4_6 (.CI(n10353), .I0(GND_net), .I1(n21_adj_1414), 
            .CO(n10354));
    SB_LUT4 i4184_4_lut (.I0(pc_data_rx[1]), .I1(r_Rx_Data), .I2(n6690), 
            .I3(n4_adj_1413), .O(n5643));   // src/uart_rx.v(49[10] 144[8])
    defparam i4184_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 led_counter_1344_1403_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_1409), .I3(n10352), .O(n127)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1344_1403_add_4_5 (.CI(n10352), .I0(GND_net), .I1(n22_adj_1409), 
            .CO(n10353));
    SB_LUT4 i4185_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[2]), .I2(n4_adj_1415), 
            .I3(n5019), .O(n5644));   // src/uart_rx.v(49[10] 144[8])
    defparam i4185_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 led_counter_1344_1403_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_1410), .I3(n10351), .O(n128)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1344_1403_add_4_4 (.CI(n10351), .I0(GND_net), .I1(n23_adj_1410), 
            .CO(n10352));
    SB_LUT4 led_counter_1344_1403_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24), .I3(n10350), .O(n129)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1344_1403_add_4_3 (.CI(n10350), .I0(GND_net), .I1(n24), 
            .CO(n10351));
    SB_LUT4 led_counter_1344_1403_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25), .I3(VCC_net), .O(n130)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1344_1403_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1344_1403_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(n25), .CO(n10350));
    SB_LUT4 i1_2_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_1401));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFF reset_clk_counter_i3_1345__i3 (.Q(reset_clk_counter[3]), .C(SLM_CLK_c), 
           .D(n10467));   // src/top.v(259[27:51])
    SB_LUT4 i4259_4_lut (.I0(\REG.mem_22_0 ), .I1(DEBUG_3_c_0), .I2(n33), 
            .I3(wr_addr_r[4]), .O(n5718));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4259_4_lut.LUT_INIT = 16'hcaaa;
    SB_DFF reset_clk_counter_i3_1345__i2 (.Q(reset_clk_counter[2]), .C(SLM_CLK_c), 
           .D(n10471));   // src/top.v(259[27:51])
    SB_DFF reset_clk_counter_i3_1345__i1 (.Q(reset_clk_counter[1]), .C(SLM_CLK_c), 
           .D(n10469));   // src/top.v(259[27:51])
    SB_LUT4 i4186_4_lut (.I0(\REG.mem_11_0 ), .I1(DEBUG_3_c_0), .I2(n26), 
            .I3(wr_addr_r[4]), .O(n5645));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4186_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i4272_4_lut (.I0(\REG.mem_28_0 ), .I1(DEBUG_3_c_0), .I2(n28), 
            .I3(wr_addr_r[4]), .O(n5731));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4272_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i12_4_lut_adj_131 (.I0(n11362), .I1(state[3]), .I2(n11257), 
            .I3(state[0]), .O(n10668));   // src/timing_controller.v(154[8] 230[4])
    defparam i12_4_lut_adj_131.LUT_INIT = 16'hcac0;
    SB_LUT4 i4189_3_lut (.I0(tx_addr_byte[7]), .I1(tx_data_byte[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5648));   // src/top.v(1165[8] 1232[4])
    defparam i4189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4190_3_lut (.I0(tx_addr_byte[6]), .I1(tx_data_byte[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5649));   // src/top.v(1165[8] 1232[4])
    defparam i4190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4191_3_lut (.I0(tx_addr_byte[5]), .I1(tx_data_byte[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5650));   // src/top.v(1165[8] 1232[4])
    defparam i4191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4192_3_lut (.I0(tx_addr_byte[4]), .I1(tx_data_byte[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5651));   // src/top.v(1165[8] 1232[4])
    defparam i4192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4193_3_lut (.I0(tx_addr_byte[3]), .I1(tx_data_byte[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5652));   // src/top.v(1165[8] 1232[4])
    defparam i4193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4194_3_lut (.I0(tx_addr_byte[2]), .I1(tx_data_byte[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5653));   // src/top.v(1165[8] 1232[4])
    defparam i4194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4195_3_lut (.I0(tx_addr_byte[1]), .I1(tx_data_byte[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5654));   // src/top.v(1165[8] 1232[4])
    defparam i4195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4196_4_lut (.I0(\REG.mem_12_0 ), .I1(DEBUG_3_c_0), .I2(n28), 
            .I3(wr_addr_r[4]), .O(n5655));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4196_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i4260_4_lut (.I0(\REG.mem_23_0 ), .I1(DEBUG_3_c_0), .I2(n35), 
            .I3(wr_addr_r[4]), .O(n5719));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4260_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i4197_4_lut (.I0(pc_data_rx[3]), .I1(r_Rx_Data), .I2(n6690), 
            .I3(n4_adj_1415), .O(n5656));   // src/uart_rx.v(49[10] 144[8])
    defparam i4197_4_lut.LUT_INIT = 16'haaca;
    GND i1 (.Y(GND_net));
    SB_LUT4 i4198_4_lut (.I0(\REG.mem_13_0 ), .I1(DEBUG_3_c_0), .I2(n30), 
            .I3(wr_addr_r[4]), .O(n5657));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4198_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i4199_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[4]), .I2(n4_adj_1407), 
            .I3(n5019), .O(n5658));   // src/uart_rx.v(49[10] 144[8])
    defparam i4199_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4200_4_lut (.I0(\REG.mem_14_0 ), .I1(DEBUG_3_c_0), .I2(n32_adj_1403), 
            .I3(wr_addr_r[4]), .O(n5659));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4200_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 reset_all_w_I_0_1_lut (.I0(reset_all_w), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(RESET_c));   // src/top.v(295[16:28])
    defparam reset_all_w_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_IO FIFO_D1_pad (.PACKAGE_PIN(FIFO_D1), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D1_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D1_pad.PULLUP = 1'b0;
    defparam FIFO_D1_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D2_pad (.PACKAGE_PIN(FIFO_D2), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D2_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D2_pad.PULLUP = 1'b0;
    defparam FIFO_D2_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D3_pad (.PACKAGE_PIN(FIFO_D3), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D3_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D3_pad.PULLUP = 1'b0;
    defparam FIFO_D3_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D4_pad (.PACKAGE_PIN(FIFO_D4), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D4_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D4_pad.PULLUP = 1'b0;
    defparam FIFO_D4_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D5_pad (.PACKAGE_PIN(FIFO_D5), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D5_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D5_pad.PULLUP = 1'b0;
    defparam FIFO_D5_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D6_pad (.PACKAGE_PIN(FIFO_D6), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D6_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D6_pad.PULLUP = 1'b0;
    defparam FIFO_D6_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D7_pad (.PACKAGE_PIN(FIFO_D7), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D7_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D7_pad.PULLUP = 1'b0;
    defparam FIFO_D7_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D8_pad (.PACKAGE_PIN(FIFO_D8), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D8_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D8_pad.PULLUP = 1'b0;
    defparam FIFO_D8_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D9_pad (.PACKAGE_PIN(FIFO_D9), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D9_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D9_pad.PULLUP = 1'b0;
    defparam FIFO_D9_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D10_pad (.PACKAGE_PIN(FIFO_D10), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D10_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D10_pad.PULLUP = 1'b0;
    defparam FIFO_D10_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D11_pad (.PACKAGE_PIN(FIFO_D11), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D11_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D11_pad.PULLUP = 1'b0;
    defparam FIFO_D11_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D12_pad (.PACKAGE_PIN(FIFO_D12), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D12_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D12_pad.PULLUP = 1'b0;
    defparam FIFO_D12_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D13_pad (.PACKAGE_PIN(FIFO_D13), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D13_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D13_pad.PULLUP = 1'b0;
    defparam FIFO_D13_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D14_pad (.PACKAGE_PIN(FIFO_D14), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D14_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D14_pad.PULLUP = 1'b0;
    defparam FIFO_D14_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D15_pad (.PACKAGE_PIN(FIFO_D15), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D15_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D15_pad.PULLUP = 1'b0;
    defparam FIFO_D15_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D15_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D16_pad (.PACKAGE_PIN(FIFO_D16), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D16_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D16_pad.PULLUP = 1'b0;
    defparam FIFO_D16_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D16_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D17_pad (.PACKAGE_PIN(FIFO_D17), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D17_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D17_pad.PULLUP = 1'b0;
    defparam FIFO_D17_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D17_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D18_pad (.PACKAGE_PIN(FIFO_D18), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D18_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D18_pad.PULLUP = 1'b0;
    defparam FIFO_D18_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D19_pad (.PACKAGE_PIN(FIFO_D19), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D19_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D19_pad.PULLUP = 1'b0;
    defparam FIFO_D19_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D20_pad (.PACKAGE_PIN(FIFO_D20), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D20_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D20_pad.PULLUP = 1'b0;
    defparam FIFO_D20_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D21_pad (.PACKAGE_PIN(FIFO_D21), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D21_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D21_pad.PULLUP = 1'b0;
    defparam FIFO_D21_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D22_pad (.PACKAGE_PIN(FIFO_D22), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D22_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D22_pad.PULLUP = 1'b0;
    defparam FIFO_D22_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D23_pad (.PACKAGE_PIN(FIFO_D23), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D23_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D23_pad.PULLUP = 1'b0;
    defparam FIFO_D23_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D24_pad (.PACKAGE_PIN(FIFO_D24), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D24_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D24_pad.PULLUP = 1'b0;
    defparam FIFO_D24_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D25_pad (.PACKAGE_PIN(FIFO_D25), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D25_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D25_pad.PULLUP = 1'b0;
    defparam FIFO_D25_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D25_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D26_pad (.PACKAGE_PIN(FIFO_D26), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D26_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D26_pad.PULLUP = 1'b0;
    defparam FIFO_D26_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D26_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO FIFO_CLK_pad (.PACKAGE_PIN(FIFO_CLK), .OUTPUT_ENABLE(VCC_net), 
            .GLOBAL_BUFFER_OUTPUT(FIFO_CLK_c));   // src/top.v(84[12:20])
    defparam FIFO_CLK_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_CLK_pad.PULLUP = 1'b0;
    defparam FIFO_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D27_pad (.PACKAGE_PIN(FIFO_D27), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D27_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D27_pad.PULLUP = 1'b0;
    defparam FIFO_D27_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D27_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D28_pad (.PACKAGE_PIN(FIFO_D28), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D28_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D28_pad.PULLUP = 1'b0;
    defparam FIFO_D28_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D28_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D29_pad (.PACKAGE_PIN(FIFO_D29), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D29_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D29_pad.PULLUP = 1'b0;
    defparam FIFO_D29_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D29_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D30_pad (.PACKAGE_PIN(FIFO_D30), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D30_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D30_pad.PULLUP = 1'b0;
    defparam FIFO_D30_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D30_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D31_pad (.PACKAGE_PIN(FIFO_D31), .OUTPUT_ENABLE(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D31_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D31_pad.PULLUP = 1'b0;
    defparam FIFO_D31_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D31_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FR_RXF_pad (.PACKAGE_PIN(FR_RXF), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FR_RXF_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FR_RXF_pad.PIN_TYPE = 6'b000001;
    defparam FR_RXF_pad.PULLUP = 1'b0;
    defparam FR_RXF_pad.NEG_TRIGGER = 1'b0;
    defparam FR_RXF_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SOUT_pad (.PACKAGE_PIN(SOUT), .OUTPUT_ENABLE(VCC_net), .D_IN_0(SOUT_c)) /* synthesis IO_FF_IN=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SOUT_pad.PIN_TYPE = 6'b000001;
    defparam SOUT_pad.PULLUP = 1'b0;
    defparam SOUT_pad.NEG_TRIGGER = 1'b0;
    defparam SOUT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UART_RX_pad (.PACKAGE_PIN(UART_RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(UART_RX_c)) /* synthesis IO_FF_IN=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UART_RX_pad.PIN_TYPE = 6'b000001;
    defparam UART_RX_pad.PULLUP = 1'b0;
    defparam UART_RX_pad.NEG_TRIGGER = 1'b0;
    defparam UART_RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_SYSCLK_pad (.PACKAGE_PIN(ICE_SYSCLK), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ICE_SYSCLK_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_SYSCLK_pad.PIN_TYPE = 6'b000001;
    defparam ICE_SYSCLK_pad.PULLUP = 1'b0;
    defparam ICE_SYSCLK_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_SYSCLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CREST_pad (.PACKAGE_PIN(ICE_CREST), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CREST_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CREST_pad.PULLUP = 1'b0;
    defparam ICE_CREST_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CREST_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CDONE_pad (.PACKAGE_PIN(ICE_CDONE), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CDONE_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CDONE_pad.PULLUP = 1'b0;
    defparam ICE_CDONE_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CDONE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CLK_pad (.PACKAGE_PIN(ICE_CLK), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CLK_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CLK_pad.PULLUP = 1'b0;
    defparam ICE_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_9_pad (.PACKAGE_PIN(DEBUG_9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_9_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_9_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_9_pad.PULLUP = 1'b0;
    defparam DEBUG_9_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_8_pad (.PACKAGE_PIN(DEBUG_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_8_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_8_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_8_pad.PULLUP = 1'b0;
    defparam DEBUG_8_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_6_pad (.PACKAGE_PIN(DEBUG_6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_6_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_6_pad.PULLUP = 1'b0;
    defparam DEBUG_6_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_5_pad (.PACKAGE_PIN(DEBUG_5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_5_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_5_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_5_pad.PULLUP = 1'b0;
    defparam DEBUG_5_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_3_pad (.PACKAGE_PIN(DEBUG_3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_3_c_0));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_3_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_3_pad.PULLUP = 1'b0;
    defparam DEBUG_3_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_2_pad (.PACKAGE_PIN(DEBUG_2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_2_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_2_pad.PULLUP = 1'b0;
    defparam DEBUG_2_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_1_pad (.PACKAGE_PIN(DEBUG_1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_1_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_1_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_1_pad.PULLUP = 1'b0;
    defparam DEBUG_1_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_0_pad (.PACKAGE_PIN(DEBUG_0), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_0_c_24));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_0_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_0_pad.PULLUP = 1'b0;
    defparam DEBUG_0_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_SIWU_pad (.PACKAGE_PIN(FT_SIWU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_SIWU_pad.PIN_TYPE = 6'b011001;
    defparam FT_SIWU_pad.PULLUP = 1'b0;
    defparam FT_SIWU_pad.NEG_TRIGGER = 1'b0;
    defparam FT_SIWU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_WR_pad (.PACKAGE_PIN(FT_WR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_WR_pad.PIN_TYPE = 6'b011001;
    defparam FT_WR_pad.PULLUP = 1'b0;
    defparam FT_WR_pad.NEG_TRIGGER = 1'b0;
    defparam FT_WR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_RD_pad (.PACKAGE_PIN(FT_RD), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(FT_RD_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_RD_pad.PIN_TYPE = 6'b011001;
    defparam FT_RD_pad.PULLUP = 1'b0;
    defparam FT_RD_pad.NEG_TRIGGER = 1'b0;
    defparam FT_RD_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_OE_pad (.PACKAGE_PIN(FT_OE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(FT_OE_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_OE_pad.PIN_TYPE = 6'b011001;
    defparam FT_OE_pad.PULLUP = 1'b0;
    defparam FT_OE_pad.NEG_TRIGGER = 1'b0;
    defparam FT_OE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA10_pad (.PACKAGE_PIN(DATA10), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA10_pad.PIN_TYPE = 6'b011001;
    defparam DATA10_pad.PULLUP = 1'b0;
    defparam DATA10_pad.NEG_TRIGGER = 1'b0;
    defparam DATA10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA9_pad (.PACKAGE_PIN(DATA9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA9_pad.PIN_TYPE = 6'b011001;
    defparam DATA9_pad.PULLUP = 1'b0;
    defparam DATA9_pad.NEG_TRIGGER = 1'b0;
    defparam DATA9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA11_pad (.PACKAGE_PIN(DATA11), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA11_pad.PIN_TYPE = 6'b011001;
    defparam DATA11_pad.PULLUP = 1'b0;
    defparam DATA11_pad.NEG_TRIGGER = 1'b0;
    defparam DATA11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA12_pad (.PACKAGE_PIN(DATA12), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA12_pad.PIN_TYPE = 6'b011001;
    defparam DATA12_pad.PULLUP = 1'b0;
    defparam DATA12_pad.NEG_TRIGGER = 1'b0;
    defparam DATA12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA13_pad (.PACKAGE_PIN(DATA13), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA13_pad.PIN_TYPE = 6'b011001;
    defparam DATA13_pad.PULLUP = 1'b0;
    defparam DATA13_pad.NEG_TRIGGER = 1'b0;
    defparam DATA13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA14_pad (.PACKAGE_PIN(DATA14), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA14_pad.PIN_TYPE = 6'b011001;
    defparam DATA14_pad.PULLUP = 1'b0;
    defparam DATA14_pad.NEG_TRIGGER = 1'b0;
    defparam DATA14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA8_pad (.PACKAGE_PIN(DATA8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA8_pad.PIN_TYPE = 6'b011001;
    defparam DATA8_pad.PULLUP = 1'b0;
    defparam DATA8_pad.NEG_TRIGGER = 1'b0;
    defparam DATA8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA15_pad (.PACKAGE_PIN(DATA15), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA15_pad.PIN_TYPE = 6'b011001;
    defparam DATA15_pad.PULLUP = 1'b0;
    defparam DATA15_pad.NEG_TRIGGER = 1'b0;
    defparam DATA15_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA16_pad (.PACKAGE_PIN(DATA16), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA16_pad.PIN_TYPE = 6'b011001;
    defparam DATA16_pad.PULLUP = 1'b0;
    defparam DATA16_pad.NEG_TRIGGER = 1'b0;
    defparam DATA16_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA7_pad (.PACKAGE_PIN(DATA7), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA7_pad.PIN_TYPE = 6'b011001;
    defparam DATA7_pad.PULLUP = 1'b0;
    defparam DATA7_pad.NEG_TRIGGER = 1'b0;
    defparam DATA7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA17_pad (.PACKAGE_PIN(DATA17), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA17_pad.PIN_TYPE = 6'b011001;
    defparam DATA17_pad.PULLUP = 1'b0;
    defparam DATA17_pad.NEG_TRIGGER = 1'b0;
    defparam DATA17_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA18_pad (.PACKAGE_PIN(DATA18), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA18_pad.PIN_TYPE = 6'b011001;
    defparam DATA18_pad.PULLUP = 1'b0;
    defparam DATA18_pad.NEG_TRIGGER = 1'b0;
    defparam DATA18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA6_pad (.PACKAGE_PIN(DATA6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA6_pad.PIN_TYPE = 6'b011001;
    defparam DATA6_pad.PULLUP = 1'b0;
    defparam DATA6_pad.NEG_TRIGGER = 1'b0;
    defparam DATA6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA19_pad (.PACKAGE_PIN(DATA19), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA19_pad.PIN_TYPE = 6'b011001;
    defparam DATA19_pad.PULLUP = 1'b0;
    defparam DATA19_pad.NEG_TRIGGER = 1'b0;
    defparam DATA19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA20_pad (.PACKAGE_PIN(DATA20), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA20_pad.PIN_TYPE = 6'b011001;
    defparam DATA20_pad.PULLUP = 1'b0;
    defparam DATA20_pad.NEG_TRIGGER = 1'b0;
    defparam DATA20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA5_pad (.PACKAGE_PIN(DATA5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA5_pad.PIN_TYPE = 6'b011001;
    defparam DATA5_pad.PULLUP = 1'b0;
    defparam DATA5_pad.NEG_TRIGGER = 1'b0;
    defparam DATA5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA21_pad (.PACKAGE_PIN(DATA21), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA21_pad.PIN_TYPE = 6'b011001;
    defparam DATA21_pad.PULLUP = 1'b0;
    defparam DATA21_pad.NEG_TRIGGER = 1'b0;
    defparam DATA21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA22_pad (.PACKAGE_PIN(DATA22), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA22_pad.PIN_TYPE = 6'b011001;
    defparam DATA22_pad.PULLUP = 1'b0;
    defparam DATA22_pad.NEG_TRIGGER = 1'b0;
    defparam DATA22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA4_pad (.PACKAGE_PIN(DATA4), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA4_pad.PIN_TYPE = 6'b011001;
    defparam DATA4_pad.PULLUP = 1'b0;
    defparam DATA4_pad.NEG_TRIGGER = 1'b0;
    defparam DATA4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA23_pad (.PACKAGE_PIN(DATA23), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA23_pad.PIN_TYPE = 6'b011001;
    defparam DATA23_pad.PULLUP = 1'b0;
    defparam DATA23_pad.NEG_TRIGGER = 1'b0;
    defparam DATA23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA24_pad (.PACKAGE_PIN(DATA24), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA24_pad.PIN_TYPE = 6'b011001;
    defparam DATA24_pad.PULLUP = 1'b0;
    defparam DATA24_pad.NEG_TRIGGER = 1'b0;
    defparam DATA24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA3_pad (.PACKAGE_PIN(DATA3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA3_pad.PIN_TYPE = 6'b011001;
    defparam DATA3_pad.PULLUP = 1'b0;
    defparam DATA3_pad.NEG_TRIGGER = 1'b0;
    defparam DATA3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA25_pad (.PACKAGE_PIN(DATA25), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA25_pad.PIN_TYPE = 6'b011001;
    defparam DATA25_pad.PULLUP = 1'b0;
    defparam DATA25_pad.NEG_TRIGGER = 1'b0;
    defparam DATA25_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA26_pad (.PACKAGE_PIN(DATA26), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA26_pad.PIN_TYPE = 6'b011001;
    defparam DATA26_pad.PULLUP = 1'b0;
    defparam DATA26_pad.NEG_TRIGGER = 1'b0;
    defparam DATA26_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA2_pad (.PACKAGE_PIN(DATA2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA2_pad.PIN_TYPE = 6'b011001;
    defparam DATA2_pad.PULLUP = 1'b0;
    defparam DATA2_pad.NEG_TRIGGER = 1'b0;
    defparam DATA2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA27_pad (.PACKAGE_PIN(DATA27), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA27_pad.PIN_TYPE = 6'b011001;
    defparam DATA27_pad.PULLUP = 1'b0;
    defparam DATA27_pad.NEG_TRIGGER = 1'b0;
    defparam DATA27_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA28_pad (.PACKAGE_PIN(DATA28), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA28_pad.PIN_TYPE = 6'b011001;
    defparam DATA28_pad.PULLUP = 1'b0;
    defparam DATA28_pad.NEG_TRIGGER = 1'b0;
    defparam DATA28_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA1_pad (.PACKAGE_PIN(DATA1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA1_pad.PIN_TYPE = 6'b011001;
    defparam DATA1_pad.PULLUP = 1'b0;
    defparam DATA1_pad.NEG_TRIGGER = 1'b0;
    defparam DATA1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA29_pad (.PACKAGE_PIN(DATA29), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA29_pad.PIN_TYPE = 6'b011001;
    defparam DATA29_pad.PULLUP = 1'b0;
    defparam DATA29_pad.NEG_TRIGGER = 1'b0;
    defparam DATA29_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA30_pad (.PACKAGE_PIN(DATA30), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA30_pad.PIN_TYPE = 6'b011001;
    defparam DATA30_pad.PULLUP = 1'b0;
    defparam DATA30_pad.NEG_TRIGGER = 1'b0;
    defparam DATA30_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA0_pad (.PACKAGE_PIN(DATA0), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA0_pad.PIN_TYPE = 6'b011001;
    defparam DATA0_pad.PULLUP = 1'b0;
    defparam DATA0_pad.NEG_TRIGGER = 1'b0;
    defparam DATA0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA31_pad (.PACKAGE_PIN(DATA31), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA31_pad.PIN_TYPE = 6'b011001;
    defparam DATA31_pad.PULLUP = 1'b0;
    defparam DATA31_pad.NEG_TRIGGER = 1'b0;
    defparam DATA31_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO VALID_pad (.PACKAGE_PIN(VALID), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VALID_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam VALID_pad.PIN_TYPE = 6'b011001;
    defparam VALID_pad.PULLUP = 1'b0;
    defparam VALID_pad.NEG_TRIGGER = 1'b0;
    defparam VALID_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SYNC_pad (.PACKAGE_PIN(SYNC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SYNC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SYNC_pad.PIN_TYPE = 6'b011001;
    defparam SYNC_pad.PULLUP = 1'b0;
    defparam SYNC_pad.NEG_TRIGGER = 1'b0;
    defparam SYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INVERT_pad (.PACKAGE_PIN(INVERT), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INVERT_c_4)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INVERT_pad.PIN_TYPE = 6'b011001;
    defparam INVERT_pad.PULLUP = 1'b0;
    defparam INVERT_pad.NEG_TRIGGER = 1'b0;
    defparam INVERT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SLM_CLK_pad (.PACKAGE_PIN(SLM_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SLM_CLK_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SLM_CLK_pad.PIN_TYPE = 6'b011001;
    defparam SLM_CLK_pad.PULLUP = 1'b0;
    defparam SLM_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam SLM_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO RESET_pad (.PACKAGE_PIN(RESET), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(RESET_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RESET_pad.PIN_TYPE = 6'b011001;
    defparam RESET_pad.PULLUP = 1'b0;
    defparam RESET_pad.NEG_TRIGGER = 1'b0;
    defparam RESET_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UPDATE_pad (.PACKAGE_PIN(UPDATE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(UPDATE_c_3));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UPDATE_pad.PIN_TYPE = 6'b011001;
    defparam UPDATE_pad.PULLUP = 1'b0;
    defparam UPDATE_pad.NEG_TRIGGER = 1'b0;
    defparam UPDATE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SDAT_pad (.PACKAGE_PIN(SDAT), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SDAT_c_15)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SDAT_pad.PIN_TYPE = 6'b011001;
    defparam SDAT_pad.PULLUP = 1'b0;
    defparam SDAT_pad.NEG_TRIGGER = 1'b0;
    defparam SDAT_pad.IO_STANDARD = "SB_LVCMOS";
=======
    SB_LUT4 i4824_3_lut (.I0(\REG.mem_21_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n12), .I3(GND_net), .O(n6298));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5511_3_lut (.I0(rx_buf_byte[4]), .I1(rx_shift_reg[4]), .I2(n3963), 
            .I3(GND_net), .O(n6985));   // src/spi.v(76[8] 221[4])
    defparam i5511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5512_3_lut (.I0(rx_buf_byte[5]), .I1(rx_shift_reg[5]), .I2(n3963), 
            .I3(GND_net), .O(n6986));   // src/spi.v(76[8] 221[4])
    defparam i5512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4825_3_lut (.I0(\REG.mem_21_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n12), .I3(GND_net), .O(n6299));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4825_3_lut.LUT_INIT = 16'hcaca;
    SB_IO UART_TX_pad (.PACKAGE_PIN(UART_TX), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(UART_TX_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UART_TX_pad.PIN_TYPE = 6'b011001;
    defparam UART_TX_pad.PULLUP = 1'b0;
    defparam UART_TX_pad.NEG_TRIGGER = 1'b0;
    defparam UART_TX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i5513_3_lut (.I0(rx_buf_byte[6]), .I1(rx_shift_reg[6]), .I2(n3963), 
            .I3(GND_net), .O(n6987));   // src/spi.v(76[8] 221[4])
    defparam i5513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4826_3_lut (.I0(\REG.mem_21_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n12), .I3(GND_net), .O(n6300));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4827_3_lut (.I0(\REG.mem_21_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n12), .I3(GND_net), .O(n6301));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4828_3_lut (.I0(\REG.mem_22_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n11), .I3(GND_net), .O(n6302));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4828_3_lut.LUT_INIT = 16'hcaca;
    SB_IO SEN_pad (.PACKAGE_PIN(SEN), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SEN_c_1)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SEN_pad.PIN_TYPE = 6'b011001;
    defparam SEN_pad.PULLUP = 1'b0;
    defparam SEN_pad.NEG_TRIGGER = 1'b0;
    defparam SEN_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4829_3_lut (.I0(\REG.mem_22_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n11), .I3(GND_net), .O(n6303));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4830_3_lut (.I0(\REG.mem_22_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n11), .I3(GND_net), .O(n6304));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5514_3_lut (.I0(rx_buf_byte[7]), .I1(rx_shift_reg[7]), .I2(n3963), 
            .I3(GND_net), .O(n6988));   // src/spi.v(76[8] 221[4])
    defparam i5514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4831_3_lut (.I0(\REG.mem_22_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n11), .I3(GND_net), .O(n6305));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5515_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n6989));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5515_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4832_3_lut (.I0(\REG.mem_22_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n11), .I3(GND_net), .O(n6306));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4833_3_lut (.I0(\REG.mem_22_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n11), .I3(GND_net), .O(n6307));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4834_3_lut (.I0(\REG.mem_22_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n11), .I3(GND_net), .O(n6308));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5516_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6990));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5516_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i12212_4_lut_4_lut (.I0(state[0]), .I1(state[2]), .I2(n12906), 
            .I3(state[1]), .O(n14242));   // src/timing_controller.v(154[8] 230[4])
    defparam i12212_4_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i4835_3_lut (.I0(\REG.mem_22_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n11), .I3(GND_net), .O(n6309));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4836_3_lut (.I0(\REG.mem_22_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n11), .I3(GND_net), .O(n6310));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4837_3_lut (.I0(\REG.mem_22_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n11), .I3(GND_net), .O(n6311));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4838_3_lut (.I0(\REG.mem_22_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n11), .I3(GND_net), .O(n6312));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5517_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n6991));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5517_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5518_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6992));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5518_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i7193_1_lut (.I0(n2075), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n8659));   // src/timing_controller.v(78[11:16])
    defparam i7193_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut (.I0(reset_clk_counter[0]), .I1(reset_clk_counter[2]), 
            .I2(reset_clk_counter[3]), .I3(reset_clk_counter[1]), .O(reset_all_w_N_61));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_1438));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1921_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n3353));   // src/top.v(1165[8] 1232[4])
    defparam i1921_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5519_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n6993));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5519_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5520_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n6994));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5520_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5521_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6995));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5521_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5522_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n6996));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5522_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5523_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6997));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5523_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5524_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n6998));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5524_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5526_2_lut (.I0(reset_per_frame), .I1(rd_addr_nxt_c_5__N_573[1]), 
            .I2(GND_net), .I3(GND_net), .O(n7000));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i5526_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4839_3_lut (.I0(\REG.mem_22_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n11), .I3(GND_net), .O(n6313));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4840_3_lut (.I0(\REG.mem_22_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n11), .I3(GND_net), .O(n6314));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5528_2_lut (.I0(reset_per_frame), .I1(rd_addr_nxt_c_5__N_573[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7002));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i5528_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4841_3_lut (.I0(\REG.mem_22_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n11), .I3(GND_net), .O(n6315));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4842_3_lut (.I0(\REG.mem_22_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n11), .I3(GND_net), .O(n6316));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4843_3_lut (.I0(\REG.mem_22_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n11), .I3(GND_net), .O(n6317));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4844_3_lut (.I0(\REG.mem_22_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n11), .I3(GND_net), .O(n6318));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5529_2_lut (.I0(reset_per_frame), .I1(rd_addr_nxt_c_5__N_573[4]), 
            .I2(GND_net), .I3(GND_net), .O(n7003));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i5529_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4845_3_lut (.I0(\REG.mem_22_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n11), .I3(GND_net), .O(n6319));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5530_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n7004));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5530_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4846_3_lut (.I0(\REG.mem_22_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n11), .I3(GND_net), .O(n6320));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4847_3_lut (.I0(\REG.mem_22_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n11), .I3(GND_net), .O(n6321));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4848_3_lut (.I0(\REG.mem_22_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n11), .I3(GND_net), .O(n6322));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4849_3_lut (.I0(\REG.mem_22_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n11), .I3(GND_net), .O(n6323));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5531_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n7005));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5531_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4850_3_lut (.I0(\REG.mem_22_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n11), .I3(GND_net), .O(n6324));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4851_3_lut (.I0(\REG.mem_22_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n11), .I3(GND_net), .O(n6325));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5532_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7006));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5532_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4852_3_lut (.I0(\REG.mem_22_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n11), .I3(GND_net), .O(n6326));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4853_3_lut (.I0(\REG.mem_22_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n11), .I3(GND_net), .O(n6327));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4853_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_addr_byte_r_i0_i7 (.Q(tx_addr_byte[7]), .C(SLM_CLK_c), .D(n7021));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_addr_byte_r_i0_i6 (.Q(tx_addr_byte[6]), .C(SLM_CLK_c), .D(n7020));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_addr_byte_r_i0_i5 (.Q(tx_addr_byte[5]), .C(SLM_CLK_c), .D(n7019));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_addr_byte_r_i0_i4 (.Q(tx_addr_byte[4]), .C(SLM_CLK_c), .D(n7018));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_addr_byte_r_i0_i3 (.Q(tx_addr_byte[3]), .C(SLM_CLK_c), .D(n7017));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_addr_byte_r_i0_i2 (.Q(tx_addr_byte[2]), .C(SLM_CLK_c), .D(n7016));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_addr_byte_r_i0_i1 (.Q(tx_addr_byte[1]), .C(SLM_CLK_c), .D(n7015));   // src/top.v(1165[8] 1232[4])
    SB_LUT4 i4854_3_lut (.I0(\REG.mem_22_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n11), .I3(GND_net), .O(n6328));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4855_3_lut (.I0(\REG.mem_22_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n11), .I3(GND_net), .O(n6329));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4856_3_lut (.I0(\REG.mem_22_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n11), .I3(GND_net), .O(n6330));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4856_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF spi_start_transfer_r_84 (.Q(spi_start_transfer_r), .C(SLM_CLK_c), 
           .D(n3468));   // src/top.v(1165[8] 1232[4])
    SB_DFF start_tx_81 (.Q(r_SM_Main_2__N_1029[0]), .C(SLM_CLK_c), .D(n6941));   // src/top.v(1001[8] 1019[4])
    SB_DFF tx_data_byte_r_i0_i1 (.Q(tx_data_byte[1]), .C(SLM_CLK_c), .D(n6938));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_data_byte_r_i0_i2 (.Q(tx_data_byte[2]), .C(SLM_CLK_c), .D(n6937));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_data_byte_r_i0_i3 (.Q(tx_data_byte[3]), .C(SLM_CLK_c), .D(n6936));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_data_byte_r_i0_i4 (.Q(tx_data_byte[4]), .C(SLM_CLK_c), .D(n6935));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_data_byte_r_i0_i5 (.Q(tx_data_byte[5]), .C(SLM_CLK_c), .D(n6934));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_data_byte_r_i0_i6 (.Q(tx_data_byte[6]), .C(SLM_CLK_c), .D(n6933));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_data_byte_r_i0_i7 (.Q(tx_data_byte[7]), .C(SLM_CLK_c), .D(n6932));   // src/top.v(1165[8] 1232[4])
    SB_LUT4 i4857_3_lut (.I0(\REG.mem_22_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n11), .I3(GND_net), .O(n6331));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4858_3_lut (.I0(\REG.mem_22_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n11), .I3(GND_net), .O(n6332));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5533_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n7007));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5533_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5534_2_lut (.I0(reset_per_frame), .I1(wr_addr_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n7008));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5534_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5446_4_lut_4_lut (.I0(rd_fifo_en_w), .I1(reset_all_w), .I2(rd_addr_p1_w_adj_1522[2]), 
            .I3(rd_addr_r_adj_1520[2]), .O(n6920));
    defparam i5446_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i5535_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n7009));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5535_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5449_4_lut_4_lut (.I0(rd_fifo_en_w), .I1(reset_all_w), .I2(rd_addr_p1_w_adj_1522[1]), 
            .I3(rd_addr_r_adj_1520[1]), .O(n6923));
    defparam i5449_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i5536_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n7010));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5536_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5537_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7011));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5537_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5538_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n7012));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5538_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5539_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n7013));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5539_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5540_2_lut (.I0(reset_per_frame_latched), .I1(n663), .I2(GND_net), 
            .I3(GND_net), .O(n7014));   // src/usb3_if.v(97[9] 199[16])
    defparam i5540_2_lut.LUT_INIT = 16'h4444;
    SB_DFF even_byte_flag_89 (.Q(even_byte_flag), .C(SLM_CLK_c), .D(n3353));   // src/top.v(1165[8] 1232[4])
    SB_LUT4 i5541_3_lut (.I0(tx_addr_byte[1]), .I1(tx_data_byte[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n7015));   // src/top.v(1165[8] 1232[4])
    defparam i5541_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5542_3_lut (.I0(tx_addr_byte[2]), .I1(tx_data_byte[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n7016));   // src/top.v(1165[8] 1232[4])
    defparam i5542_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5543_3_lut (.I0(tx_addr_byte[3]), .I1(tx_data_byte[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n7017));   // src/top.v(1165[8] 1232[4])
    defparam i5543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5544_3_lut (.I0(tx_addr_byte[4]), .I1(tx_data_byte[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n7018));   // src/top.v(1165[8] 1232[4])
    defparam i5544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5545_3_lut (.I0(tx_addr_byte[5]), .I1(tx_data_byte[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n7019));   // src/top.v(1165[8] 1232[4])
    defparam i5545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5546_3_lut (.I0(tx_addr_byte[6]), .I1(tx_data_byte[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n7020));   // src/top.v(1165[8] 1232[4])
    defparam i5546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5547_3_lut (.I0(tx_addr_byte[7]), .I1(tx_data_byte[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n7021));   // src/top.v(1165[8] 1232[4])
    defparam i5547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4859_3_lut (.I0(\REG.mem_22_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n11), .I3(GND_net), .O(n6333));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4860_3_lut (.I0(\REG.mem_23_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n10), .I3(GND_net), .O(n6334));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4861_3_lut (.I0(\REG.mem_23_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n10), .I3(GND_net), .O(n6335));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4862_3_lut (.I0(\REG.mem_23_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n10), .I3(GND_net), .O(n6336));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4862_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1434_1494__i0 (.Q(n25_adj_1437), .C(SLM_CLK_c), .D(n130));   // src/top.v(203[20:35])
    SB_LUT4 i4863_3_lut (.I0(\REG.mem_23_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n10), .I3(GND_net), .O(n6337));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4864_3_lut (.I0(\REG.mem_23_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n10), .I3(GND_net), .O(n6338));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4865_3_lut (.I0(\REG.mem_23_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n10), .I3(GND_net), .O(n6339));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4866_3_lut (.I0(\REG.mem_23_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n10), .I3(GND_net), .O(n6340));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4866_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_clk_counter_i3_1435__i0 (.Q(reset_clk_counter[0]), .C(SLM_CLK_c), 
           .D(n25_adj_1438));   // src/top.v(259[27:51])
    SB_LUT4 i4867_3_lut (.I0(\REG.mem_23_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n10), .I3(GND_net), .O(n6341));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4868_3_lut (.I0(\REG.mem_23_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n10), .I3(GND_net), .O(n6342));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4869_3_lut (.I0(\REG.mem_23_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n10), .I3(GND_net), .O(n6343));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4870_3_lut (.I0(\REG.mem_23_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n10), .I3(GND_net), .O(n6344));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4871_3_lut (.I0(\REG.mem_23_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n10), .I3(GND_net), .O(n6345));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4872_3_lut (.I0(\REG.mem_23_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n10), .I3(GND_net), .O(n6346));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4873_3_lut (.I0(\REG.mem_23_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n10), .I3(GND_net), .O(n6347));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4874_3_lut (.I0(\REG.mem_23_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n10), .I3(GND_net), .O(n6348));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4875_3_lut (.I0(\REG.mem_23_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n10), .I3(GND_net), .O(n6349));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4876_3_lut (.I0(\REG.mem_23_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n10), .I3(GND_net), .O(n6350));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4877_3_lut (.I0(\REG.mem_23_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n10), .I3(GND_net), .O(n6351));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4878_3_lut (.I0(\REG.mem_23_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n10), .I3(GND_net), .O(n6352));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4879_3_lut (.I0(\REG.mem_23_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n10), .I3(GND_net), .O(n6353));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4880_3_lut (.I0(\REG.mem_23_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n10), .I3(GND_net), .O(n6354));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4881_3_lut (.I0(\REG.mem_23_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n10), .I3(GND_net), .O(n6355));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4882_3_lut (.I0(\REG.mem_23_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n10), .I3(GND_net), .O(n6356));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4883_3_lut (.I0(\REG.mem_23_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n10), .I3(GND_net), .O(n6357));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4884_3_lut (.I0(\REG.mem_23_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n10), .I3(GND_net), .O(n6358));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4885_3_lut (.I0(\REG.mem_23_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n10), .I3(GND_net), .O(n6359));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4886_3_lut (.I0(\REG.mem_23_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n10), .I3(GND_net), .O(n6360));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4887_3_lut (.I0(\REG.mem_23_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n10), .I3(GND_net), .O(n6361));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4888_3_lut (.I0(\REG.mem_23_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n10), .I3(GND_net), .O(n6362));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4889_3_lut (.I0(\REG.mem_23_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n10), .I3(GND_net), .O(n6363));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4890_3_lut (.I0(\REG.mem_23_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n10), .I3(GND_net), .O(n6364));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4891_3_lut (.I0(\REG.mem_23_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n10), .I3(GND_net), .O(n6365));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4892_3_lut (.I0(\REG.mem_24_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n9), .I3(GND_net), .O(n6366));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4893_3_lut (.I0(\REG.mem_24_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n9), .I3(GND_net), .O(n6367));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4894_3_lut (.I0(\REG.mem_24_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n9), .I3(GND_net), .O(n6368));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4895_3_lut (.I0(\REG.mem_24_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n9), .I3(GND_net), .O(n6369));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4896_3_lut (.I0(\REG.mem_24_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n9), .I3(GND_net), .O(n6370));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4897_3_lut (.I0(\REG.mem_24_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n9), .I3(GND_net), .O(n6371));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4898_3_lut (.I0(\REG.mem_24_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n9), .I3(GND_net), .O(n6372));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4899_3_lut (.I0(\REG.mem_24_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n9), .I3(GND_net), .O(n6373));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4900_3_lut (.I0(\REG.mem_24_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n9), .I3(GND_net), .O(n6374));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4901_3_lut (.I0(\REG.mem_24_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n9), .I3(GND_net), .O(n6375));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4902_3_lut (.I0(\REG.mem_24_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n9), .I3(GND_net), .O(n6376));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4903_3_lut (.I0(\REG.mem_24_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n9), .I3(GND_net), .O(n6377));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4904_3_lut (.I0(\REG.mem_24_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n9), .I3(GND_net), .O(n6378));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4905_3_lut (.I0(\REG.mem_24_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n9), .I3(GND_net), .O(n6379));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4906_3_lut (.I0(\REG.mem_24_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n9), .I3(GND_net), .O(n6380));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4907_3_lut (.I0(\REG.mem_24_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n9), .I3(GND_net), .O(n6381));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4908_3_lut (.I0(\REG.mem_24_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n9), .I3(GND_net), .O(n6382));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4909_3_lut (.I0(\REG.mem_24_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n9), .I3(GND_net), .O(n6383));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1434_1494_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(DEBUG_0_c_24), .I3(n12177), .O(n106)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 led_counter_1434_1494_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n2), .I3(n12176), .O(n107)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_25 (.CI(n12176), .I0(GND_net), 
            .I1(n2), .CO(n12177));
    SB_LUT4 led_counter_1434_1494_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3), .I3(n12175), .O(n108)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_24_lut.LUT_INIT = 16'hC33C;
>>>>>>> Stashed changes
    SB_IO SCK_pad (.PACKAGE_PIN(SCK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SCK_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SCK_pad.PIN_TYPE = 6'b011001;
    defparam SCK_pad.PULLUP = 1'b0;
    defparam SCK_pad.NEG_TRIGGER = 1'b0;
    defparam SCK_pad.IO_STANDARD = "SB_LVCMOS";
<<<<<<< Updated upstream
    SB_IO SEN_pad (.PACKAGE_PIN(SEN), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SEN_c_1)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SEN_pad.PIN_TYPE = 6'b011001;
    defparam SEN_pad.PULLUP = 1'b0;
    defparam SEN_pad.NEG_TRIGGER = 1'b0;
    defparam SEN_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4202_4_lut (.I0(\REG.mem_15_0 ), .I1(DEBUG_3_c_0), .I2(n34), 
            .I3(wr_addr_r[4]), .O(n5661));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4202_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i4203_4_lut (.I0(\REG.mem_16_0 ), .I1(DEBUG_3_c_0), .I2(n21), 
            .I3(wr_addr_r[4]), .O(n5662));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4203_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i4204_2_lut (.I0(reset_per_frame), .I1(wr_grey_w[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5663));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    defparam i4204_2_lut.LUT_INIT = 16'h4444;
    SB_DFF tx_addr_byte_r_i0_i1 (.Q(tx_addr_byte[1]), .C(SLM_CLK_c), .D(n5654));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_addr_byte_r_i0_i2 (.Q(tx_addr_byte[2]), .C(SLM_CLK_c), .D(n5653));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_addr_byte_r_i0_i3 (.Q(tx_addr_byte[3]), .C(SLM_CLK_c), .D(n5652));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_addr_byte_r_i0_i4 (.Q(tx_addr_byte[4]), .C(SLM_CLK_c), .D(n5651));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_addr_byte_r_i0_i5 (.Q(tx_addr_byte[5]), .C(SLM_CLK_c), .D(n5650));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_addr_byte_r_i0_i6 (.Q(tx_addr_byte[6]), .C(SLM_CLK_c), .D(n5649));   // src/top.v(1165[8] 1232[4])
    SB_LUT4 i4205_4_lut (.I0(\REG.mem_17_0 ), .I1(DEBUG_3_c_0), .I2(n23_adj_1402), 
            .I3(wr_addr_r[4]), .O(n5664));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4205_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i4261_3_lut (.I0(tx_data_byte[3]), .I1(pc_data_rx[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5720));   // src/top.v(1165[8] 1232[4])
    defparam i4261_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_addr_byte_r_i0_i7 (.Q(tx_addr_byte[7]), .C(SLM_CLK_c), .D(n5648));   // src/top.v(1165[8] 1232[4])
    SB_LUT4 i4206_4_lut (.I0(pc_data_rx[5]), .I1(r_Rx_Data), .I2(n6690), 
            .I3(n4_adj_1407), .O(n5665));   // src/uart_rx.v(49[10] 144[8])
    defparam i4206_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i4207_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5666));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4207_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4208_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5667));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4208_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4209_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5668));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4209_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4210_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5669));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4210_2_lut.LUT_INIT = 16'h4444;
    SB_DFF reset_clk_counter_i3_1345__i0 (.Q(reset_clk_counter[0]), .C(SLM_CLK_c), 
           .D(n25_adj_1401));   // src/top.v(259[27:51])
    SB_LUT4 i4211_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5670));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4211_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8779_2_lut_3_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(reset_clk_counter[1]), .I3(GND_net), .O(n10209));   // src/top.v(259[27:51])
    defparam i8779_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(reset_clk_counter[1]), .I3(GND_net), .O(n10469));   // src/top.v(259[27:51])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 i4165_2_lut_4_lut (.I0(reset_per_frame), .I1(rd_addr_r[0]), 
            .I2(rd_addr_p1_w[0]), .I3(rd_fifo_en_w), .O(n5624));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i4165_2_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4282_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[3]), 
            .I2(\mem_LUT.data_raw_r [3]), .I3(n5159), .O(n5741));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4282_4_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4286_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[4]), 
            .I2(\mem_LUT.data_raw_r [4]), .I3(n5159), .O(n5745));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4286_4_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4289_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[5]), 
            .I2(\mem_LUT.data_raw_r [5]), .I3(n5159), .O(n5748));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4289_4_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4212_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5671));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4212_2_lut.LUT_INIT = 16'h4444;
    SB_DFF led_counter_1344_1403__i24 (.Q(DEBUG_0_c_24), .C(SLM_CLK_c), 
           .D(n106_adj_1406));   // src/top.v(203[20:35])
    SB_LUT4 i4262_4_lut (.I0(\REG.mem_24_0 ), .I1(DEBUG_3_c_0), .I2(n20), 
            .I3(wr_addr_r[4]), .O(n5721));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4262_4_lut.LUT_INIT = 16'hcaaa;
    SB_DFF spi_start_transfer_r_84 (.Q(spi_start_transfer_r), .C(SLM_CLK_c), 
           .D(n3426));   // src/top.v(1165[8] 1232[4])
    SB_LUT4 i4213_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5672));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4213_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4214_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5673));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4214_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4353_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[0]), 
            .I2(\mem_LUT.data_raw_r [0]), .I3(n5159), .O(n5812));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4353_4_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4215_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5674));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4215_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut (.I0(reset_clk_counter[2]), .I1(reset_all_w_N_61), 
            .I2(reset_clk_counter[0]), .I3(reset_clk_counter[1]), .O(n10471));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'haaa6;
    SB_LUT4 i4158_4_lut_4_lut (.I0(tx_uart_active_flag), .I1(r_SM_Main_adj_1435[1]), 
            .I2(r_SM_Main_adj_1435[2]), .I3(n11079), .O(n5617));   // src/uart_tx.v(38[10] 141[8])
    defparam i4158_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i4296_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[6]), 
            .I2(\mem_LUT.data_raw_r [6]), .I3(n5159), .O(n5755));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4296_4_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4349_3_lut_4_lut (.I0(r_SM_Main_2__N_1028[0]), .I1(fifo_read_cmd), 
            .I2(is_fifo_empty_flag), .I3(tx_uart_active_flag), .O(n5808));   // src/top.v(1001[8] 1019[4])
    defparam i4349_3_lut_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4302_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[7]), 
            .I2(\mem_LUT.data_raw_r [7]), .I3(n5159), .O(n5761));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4302_4_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4264_4_lut (.I0(\REG.mem_25_0 ), .I1(DEBUG_3_c_0), .I2(n22), 
            .I3(wr_addr_r[4]), .O(n5723));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4264_4_lut.LUT_INIT = 16'hcaaa;
    SB_DFF led_counter_1344_1403__i23 (.Q(n2), .C(SLM_CLK_c), .D(n107));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i22 (.Q(n3_adj_1411), .C(SLM_CLK_c), .D(n108));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i21 (.Q(n4_adj_1418), .C(SLM_CLK_c), .D(n109));   // src/top.v(203[20:35])
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(rd_fifo_en_prev_r), .I1(fifo_read_cmd), 
            .I2(is_fifo_empty_flag), .I3(reset_all_w), .O(n5159));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hffae;
    SB_DFF led_counter_1344_1403__i20 (.Q(n5), .C(SLM_CLK_c), .D(n110));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i19 (.Q(n6_adj_1408), .C(SLM_CLK_c), .D(n111));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i18 (.Q(n7_adj_1412), .C(SLM_CLK_c), .D(n112));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i17 (.Q(n8), .C(SLM_CLK_c), .D(n113));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i16 (.Q(n9), .C(SLM_CLK_c), .D(n114));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i15 (.Q(n10), .C(SLM_CLK_c), .D(n115));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i14 (.Q(n11), .C(SLM_CLK_c), .D(n116));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i13 (.Q(n12), .C(SLM_CLK_c), .D(n117));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i12 (.Q(n13), .C(SLM_CLK_c), .D(n118));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i11 (.Q(n14), .C(SLM_CLK_c), .D(n119));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i10 (.Q(n15_adj_1417), .C(SLM_CLK_c), 
           .D(n120));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i9 (.Q(n16), .C(SLM_CLK_c), .D(n121));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i8 (.Q(n17), .C(SLM_CLK_c), .D(n122));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i7 (.Q(n18), .C(SLM_CLK_c), .D(n123));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i6 (.Q(n19), .C(SLM_CLK_c), .D(n124));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i5 (.Q(n20_adj_1416), .C(SLM_CLK_c), .D(n125));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i4 (.Q(n21_adj_1414), .C(SLM_CLK_c), .D(n126));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i3 (.Q(n22_adj_1409), .C(SLM_CLK_c), .D(n127));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i2 (.Q(n23_adj_1410), .C(SLM_CLK_c), .D(n128));   // src/top.v(203[20:35])
    SB_DFF led_counter_1344_1403__i1 (.Q(n24), .C(SLM_CLK_c), .D(n129));   // src/top.v(203[20:35])
    SB_LUT4 i4216_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5675));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4216_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3_4_lut (.I0(reset_clk_counter[0]), .I1(reset_clk_counter[2]), 
            .I2(reset_clk_counter[3]), .I3(reset_clk_counter[1]), .O(reset_all_w_N_61));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4265_3_lut (.I0(tx_data_byte[2]), .I1(pc_data_rx[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5724));   // src/top.v(1165[8] 1232[4])
    defparam i4265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4151_4_lut_4_lut (.I0(reset_all_w), .I1(rd_addr_r_adj_1493[1]), 
            .I2(rd_addr_r_adj_1493[0]), .I3(empty_o_N_1333), .O(n5610));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i4151_4_lut_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i1_3_lut_adj_132 (.I0(n63), .I1(state[3]), .I2(n4943), .I3(GND_net), 
            .O(n1967));   // src/timing_controller.v(78[11:16])
    defparam i1_3_lut_adj_132.LUT_INIT = 16'h2828;
    SB_DFF fifo_write_cmd_79 (.Q(fifo_write_cmd), .C(SLM_CLK_c), .D(n5632));   // src/top.v(980[8] 989[4])
    SB_LUT4 i4276_4_lut (.I0(\REG.mem_29_0 ), .I1(DEBUG_3_c_0), .I2(n30), 
            .I3(wr_addr_r[4]), .O(n5735));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4276_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i4266_4_lut (.I0(\REG.mem_26_0 ), .I1(DEBUG_3_c_0), .I2(n24_adj_1404), 
            .I3(wr_addr_r[4]), .O(n5725));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4266_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i9617_2_lut (.I0(tx_data_byte[5]), .I1(tx_data_byte[7]), .I2(GND_net), 
            .I3(GND_net), .O(n11193));
    defparam i9617_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i9683_4_lut (.I0(tx_data_byte[3]), .I1(tx_data_byte[2]), .I2(tx_data_byte[4]), 
            .I3(n11193), .O(n11261));
    defparam i9683_4_lut.LUT_INIT = 16'h8000;
    SB_DFF tx_addr_byte_r_i0_i0 (.Q(tx_addr_byte[0]), .C(SLM_CLK_c), .D(n5628));   // src/top.v(1165[8] 1232[4])
    SB_LUT4 i9940_4_lut (.I0(tx_data_byte[0]), .I1(tx_data_byte[1]), .I2(tx_data_byte[6]), 
            .I3(n11261), .O(multi_byte_spi_trans_flag_r_N_72));   // src/top.v(1214[10:31])
    defparam i9940_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i4283_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5742));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4283_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4290_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5749));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4290_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4291_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5750));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4291_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4292_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5751));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4292_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_133 (.I0(n63), .I1(n23), .I2(n4943), .I3(state[3]), 
            .O(n2072));   // src/timing_controller.v(78[11:16])
    defparam i1_4_lut_adj_133.LUT_INIT = 16'h0544;
    SB_DFF uart_rx_complete_rising_edge_82 (.Q(uart_rx_complete_rising_edge), 
           .C(SLM_CLK_c), .D(n5620));   // src/top.v(1156[8] 1162[4])
    SB_DFF start_tx_81 (.Q(r_SM_Main_2__N_1028[0]), .C(SLM_CLK_c), .D(n5808));   // src/top.v(1001[8] 1019[4])
    SB_LUT4 i4293_3_lut (.I0(tx_data_byte[7]), .I1(pc_data_rx[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5752));   // src/top.v(1165[8] 1232[4])
    defparam i4293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4218_2_lut (.I0(reset_per_frame), .I1(rd_addr_nxt_c_5__N_572[4]), 
            .I2(GND_net), .I3(GND_net), .O(n5677));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i4218_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_3_lut_adj_134 (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(reset_all_w), .I3(GND_net), .O(empty_o_N_1333));
    defparam i1_2_lut_3_lut_adj_134.LUT_INIT = 16'hf2f2;
    SB_LUT4 i4220_2_lut (.I0(reset_per_frame), .I1(rd_addr_nxt_c_5__N_572[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5679));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i4220_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3998_1_lut_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n5457));   // src/top.v(1165[8] 1232[4])
    defparam i3998_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_DFF led_counter_1344_1403__i0 (.Q(n25), .C(SLM_CLK_c), .D(n130));   // src/top.v(203[20:35])
    SB_LUT4 i4297_3_lut (.I0(tx_data_byte[6]), .I1(pc_data_rx[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5756));   // src/top.v(1165[8] 1232[4])
    defparam i4297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4298_3_lut (.I0(tx_data_byte[5]), .I1(pc_data_rx[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5757));   // src/top.v(1165[8] 1232[4])
    defparam i4298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4299_3_lut (.I0(tx_data_byte[4]), .I1(pc_data_rx[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5758));   // src/top.v(1165[8] 1232[4])
    defparam i4299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4146_3_lut (.I0(tx_data_byte[0]), .I1(pc_data_rx[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5605));   // src/top.v(1165[8] 1232[4])
    defparam i4146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4303_4_lut (.I0(\REG.mem_30_0 ), .I1(DEBUG_3_c_0), .I2(n32_adj_1403), 
            .I3(wr_addr_r[4]), .O(n5762));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4303_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i4148_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5607));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4148_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4307_4_lut (.I0(\REG.mem_31_0 ), .I1(DEBUG_3_c_0), .I2(n34), 
            .I3(wr_addr_r[4]), .O(n5766));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4307_4_lut.LUT_INIT = 16'hcaaa;
    SB_DFF tx_data_byte_r_i0_i0 (.Q(tx_data_byte[0]), .C(SLM_CLK_c), .D(n5605));   // src/top.v(1165[8] 1232[4])
    SB_LUT4 i3_4_lut_adj_135 (.I0(n63), .I1(state[1]), .I2(state[2]), 
            .I3(n11101), .O(n11700));   // src/timing_controller.v(160[5] 229[12])
    defparam i3_4_lut_adj_135.LUT_INIT = 16'h0400;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_1435[2]), .I1(r_SM_Main_2__N_1025[1]), 
            .I2(r_SM_Main_adj_1435[0]), .I3(r_SM_Main_adj_1435[1]), .O(n11691));   // src/uart_tx.v(38[10] 141[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h4000;
    SB_DFF tx_data_byte_r_i0_i4 (.Q(tx_data_byte[4]), .C(SLM_CLK_c), .D(n5758));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_data_byte_r_i0_i5 (.Q(tx_data_byte[5]), .C(SLM_CLK_c), .D(n5757));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_data_byte_r_i0_i6 (.Q(tx_data_byte[6]), .C(SLM_CLK_c), .D(n5756));   // src/top.v(1165[8] 1232[4])
    SB_DFF tx_data_byte_r_i0_i7 (.Q(tx_data_byte[7]), .C(SLM_CLK_c), .D(n5752));   // src/top.v(1165[8] 1232[4])
    SB_LUT4 i4155_4_lut (.I0(RESET_c), .I1(rd_addr_r_adj_1493[2]), .I2(rd_addr_p1_w_adj_1495[2]), 
            .I3(empty_o_N_1333), .O(n5614));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i4155_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i4267_4_lut (.I0(\REG.mem_27_0 ), .I1(DEBUG_3_c_0), .I2(n26), 
            .I3(wr_addr_r[4]), .O(n5726));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4267_4_lut.LUT_INIT = 16'hcaaa;
    \uart_rx(CLKS_PER_BIT=20)  pc_rx (.SLM_CLK_c(SLM_CLK_c), .r_SM_Main({r_SM_Main}), 
            .\r_SM_Main_2__N_949[2] (r_SM_Main_2__N_949[2]), .GND_net(GND_net), 
            .n8012(n8012), .r_Rx_Data(r_Rx_Data), .n5214(n5214), .n4(n4_adj_1413), 
            .n5709(n5709), .pc_data_rx({pc_data_rx}), .n5692(n5692), .n5527(n5527), 
            .n4_adj_1(n4_adj_1415), .UART_RX_c(UART_RX_c), .n5665(n5665), 
            .n5658(n5658), .n5656(n5656), .n4_adj_2(n4_adj_1407), .\r_Bit_Index[0] (r_Bit_Index[0]), 
            .n6690(n6690), .n5644(n5644), .n5643(n5643), .n5825(n5825), 
            .n10608(n10608), .VCC_net(VCC_net), .debug_led3(debug_led3), 
            .n5821(n5821), .n5019(n5019)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(790[42] 795[3])
    SB_LUT4 i4271_3_lut (.I0(tx_data_byte[1]), .I1(pc_data_rx[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5730));   // src/top.v(1165[8] 1232[4])
    defparam i4271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9863_2_lut_3_lut (.I0(state[2]), .I1(state[3]), .I2(state[1]), 
            .I3(GND_net), .O(n11362));   // src/timing_controller.v(154[8] 230[4])
    defparam i9863_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFFSR multi_byte_spi_trans_flag_r_86 (.Q(multi_byte_spi_trans_flag_r), 
            .C(SLM_CLK_c), .D(multi_byte_spi_trans_flag_r_N_72), .R(n5457));   // src/top.v(1165[8] 1232[4])
    SB_LUT4 i4222_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5681));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4222_2_lut.LUT_INIT = 16'h4444;
    clock clock_inst (.GND_net(GND_net), .VCC_net(VCC_net), .ICE_SYSCLK_c(ICE_SYSCLK_c), 
          .pll_clk_unbuf(pll_clk_unbuf)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(222[7] 228[3])
    SB_LUT4 i4275_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[1]), 
            .I2(\mem_LUT.data_raw_r [1]), .I3(n5159), .O(n5734));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4275_4_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i1_4_lut_4_lut (.I0(is_tx_fifo_full_flag), .I1(n11239), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h2222;
    SB_DFF fifo_read_cmd_80 (.Q(fifo_read_cmd), .C(SLM_CLK_c), .D(start_tx_N_64));   // src/top.v(1001[8] 1019[4])
    SB_LUT4 i4223_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5682));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4223_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_949[2]), 
            .I3(r_SM_Main[0]), .O(n5101));   // src/uart_rx.v(49[10] 144[8])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i4224_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5683));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4224_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1376_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(reset_all_w), .I3(GND_net), .O(n2704));
    defparam i1376_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i6611_2_lut_3_lut (.I0(state[1]), .I1(state[0]), .I2(n63), 
            .I3(GND_net), .O(n8057));
    defparam i6611_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i4225_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5684));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4225_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i39_3_lut_4_lut_3_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(GND_net), .O(n23));
    defparam i39_3_lut_4_lut_3_lut.LUT_INIT = 16'h8686;
    SB_LUT4 i4310_4_lut (.I0(RESET_c), .I1(wr_addr_r_adj_1490[2]), .I2(wr_addr_p1_w_adj_1492[2]), 
            .I3(n2704), .O(n5769));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i4310_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i4226_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5685));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4226_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4279_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[2]), 
            .I2(\mem_LUT.data_raw_r [2]), .I3(n5159), .O(n5738));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4279_4_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4227_4_lut (.I0(\REG.mem_18_0 ), .I1(DEBUG_3_c_0), .I2(n25_adj_1405), 
            .I3(wr_addr_r[4]), .O(n5686));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4227_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i4228_2_lut (.I0(reset_per_frame), .I1(rd_addr_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5687));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4228_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4229_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5688));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4229_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4174_2_lut_3_lut (.I0(reset_all_w), .I1(fifo_read_cmd), .I2(is_fifo_empty_flag), 
            .I3(GND_net), .O(n5633));   // src/fifo_quad_word_mod.v(353[29] 363[32])
    defparam i4174_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i4230_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5689));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4230_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4231_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5690));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4231_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i9937_2_lut (.I0(is_fifo_empty_flag), .I1(tx_uart_active_flag), 
            .I2(GND_net), .I3(GND_net), .O(start_tx_N_64));
    defparam i9937_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i4232_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5691));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4232_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4152_4_lut (.I0(\REG.mem_0_0 ), .I1(DEBUG_3_c_0), .I2(n21), 
            .I3(wr_addr_r[4]), .O(n5611));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4152_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i4156_4_lut (.I0(\REG.mem_2_0 ), .I1(DEBUG_3_c_0), .I2(n25_adj_1405), 
            .I3(wr_addr_r[4]), .O(n5615));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4156_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i4157_2_lut (.I0(bluejay_data_out_31__N_919), .I1(bluejay_data_out_31__N_920), 
            .I2(GND_net), .I3(GND_net), .O(n5616));   // src/bluejay_data.v(134[8] 156[4])
    defparam i4157_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6394_1_lut (.I0(n1967), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n7836));   // src/timing_controller.v(78[11:16])
    defparam i6394_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4159_3_lut (.I0(r_Tx_Data[0]), .I1(fifo_temp_output[0]), .I2(n4715), 
            .I3(GND_net), .O(n5618));   // src/uart_tx.v(38[10] 141[8])
    defparam i4159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4233_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[6]), .I2(n8012), 
            .I3(n5019), .O(n5692));   // src/uart_rx.v(49[10] 144[8])
    defparam i4233_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i4161_2_lut (.I0(uart_rx_complete_prev), .I1(debug_led3), .I2(GND_net), 
            .I3(GND_net), .O(n5620));   // src/top.v(1156[8] 1162[4])
    defparam i4161_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4234_3_lut (.I0(rx_buf_byte[7]), .I1(rx_shift_reg[7]), .I2(n5120), 
            .I3(GND_net), .O(n5693));   // src/spi.v(76[8] 221[4])
    defparam i4234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4162_3_lut (.I0(rx_buf_byte[0]), .I1(rx_shift_reg[0]), .I2(n5120), 
            .I3(GND_net), .O(n5621));   // src/spi.v(76[8] 221[4])
    defparam i4162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4163_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5622));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4163_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4235_3_lut (.I0(rx_buf_byte[6]), .I1(rx_shift_reg[6]), .I2(n5120), 
            .I3(GND_net), .O(n5694));   // src/spi.v(76[8] 221[4])
    defparam i4235_3_lut.LUT_INIT = 16'hcaca;
    spi spi0 (.VCC_net(VCC_net), .GND_net(GND_net), .SLM_CLK_c(SLM_CLK_c), 
        .SEN_c_1(SEN_c_1), .SOUT_c(SOUT_c), .n5113(n5113), .\rx_shift_reg[0] (rx_shift_reg[0]), 
        .n2329(n2329), .multi_byte_spi_trans_flag_r(multi_byte_spi_trans_flag_r), 
        .spi_start_transfer_r(spi_start_transfer_r), .tx_addr_byte({tx_addr_byte}), 
        .n5081(n5081), .SDAT_c_15(SDAT_c_15), .n5706(n5706), .\rx_shift_reg[1] (rx_shift_reg[1]), 
        .n5705(n5705), .\rx_shift_reg[2] (rx_shift_reg[2]), .n5704(n5704), 
        .\rx_shift_reg[3] (rx_shift_reg[3]), .n5703(n5703), .\rx_shift_reg[4] (rx_shift_reg[4]), 
        .n5702(n5702), .\rx_shift_reg[5] (rx_shift_reg[5]), .n5701(n5701), 
        .\rx_shift_reg[6] (rx_shift_reg[6]), .n5700(n5700), .\rx_shift_reg[7] (rx_shift_reg[7]), 
        .n5699(n5699), .rx_buf_byte({rx_buf_byte}), .n5698(n5698), .n5697(n5697), 
        .n5696(n5696), .n5695(n5695), .n5694(n5694), .\tx_data_byte[1] (tx_data_byte[1]), 
        .\tx_shift_reg[0] (tx_shift_reg[0]), .\tx_data_byte[2] (tx_data_byte[2]), 
        .\tx_data_byte[3] (tx_data_byte[3]), .\tx_data_byte[4] (tx_data_byte[4]), 
        .n5693(n5693), .\tx_data_byte[5] (tx_data_byte[5]), .\tx_data_byte[6] (tx_data_byte[6]), 
        .\tx_data_byte[7] (tx_data_byte[7]), .spi_rx_byte_ready(spi_rx_byte_ready), 
        .SCK_c_0(SCK_c_0), .n5120(n5120), .n10792(n10792), .n5621(n5621)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(924[5] 948[2])
    usb3_if usb3_if_inst (.reset_per_frame(reset_per_frame), .SLM_CLK_c(SLM_CLK_c), 
            .DEBUG_9_c(DEBUG_9_c), .VCC_net(VCC_net), .FT_RD_c(FT_RD_c), 
            .FIFO_CLK_c(FIFO_CLK_c), .DEBUG_3_c_0(DEBUG_3_c_0), .dc32_fifo_write_enable(dc32_fifo_write_enable), 
            .buffer_switch_done(buffer_switch_done), .buffer_switch_done_latched(buffer_switch_done_latched), 
            .FT_OE_c(FT_OE_c), .FR_RXF_c(FR_RXF_c), .GND_net(GND_net), 
            .DEBUG_1_c(DEBUG_1_c), .FIFO_D0_c_0(FIFO_D0_c_0)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(544[9] 560[3])
    fifo_sc_32_lut_gen fifo_sc_32_lut_gen_inst (.SLM_CLK_c(SLM_CLK_c), .sc32_fifo_almost_empty(sc32_fifo_almost_empty), 
            .reset_all(reset_all), .GND_net(GND_net), .dc32_fifo_read_enable(dc32_fifo_read_enable), 
            .sc32_fifo_read_enable(sc32_fifo_read_enable)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(620[20] 634[2])
    SB_LUT4 i1_3_lut_adj_136 (.I0(reset_clk_counter[3]), .I1(reset_clk_counter[2]), 
            .I2(n10209), .I3(GND_net), .O(n10467));
    defparam i1_3_lut_adj_136.LUT_INIT = 16'ha9a9;
    SB_LUT4 i4236_3_lut (.I0(rx_buf_byte[5]), .I1(rx_shift_reg[5]), .I2(n5120), 
            .I3(GND_net), .O(n5695));   // src/spi.v(76[8] 221[4])
    defparam i4236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4237_3_lut (.I0(rx_buf_byte[4]), .I1(rx_shift_reg[4]), .I2(n5120), 
            .I3(GND_net), .O(n5696));   // src/spi.v(76[8] 221[4])
    defparam i4237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4358_3_lut (.I0(n5525), .I1(r_Bit_Index_adj_1437[0]), .I2(n5212), 
            .I3(GND_net), .O(n5817));   // src/uart_tx.v(38[10] 141[8])
    defparam i4358_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i4238_3_lut (.I0(rx_buf_byte[3]), .I1(rx_shift_reg[3]), .I2(n5120), 
            .I3(GND_net), .O(n5697));   // src/spi.v(76[8] 221[4])
    defparam i4238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4239_3_lut (.I0(rx_buf_byte[2]), .I1(rx_shift_reg[2]), .I2(n5120), 
            .I3(GND_net), .O(n5698));   // src/spi.v(76[8] 221[4])
    defparam i4239_3_lut.LUT_INIT = 16'hcaca;
    FIFO_Quad_Word tx_fifo (.rd_addr_r({rd_addr_r_adj_1493}), .SLM_CLK_c(SLM_CLK_c), 
            .reset_all_w(reset_all_w), .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r [0]), 
            .wr_addr_r({wr_addr_r_adj_1490}), .fifo_write_cmd(fifo_write_cmd), 
            .is_tx_fifo_full_flag(is_tx_fifo_full_flag), .wr_fifo_en_w(wr_fifo_en_w), 
            .GND_net(GND_net), .n2704(n2704), .\wr_addr_p1_w[2] (wr_addr_p1_w_adj_1492[2]), 
            .n1(n1), .n10381(n10381), .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r [7]), 
            .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r [6]), .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r [5]), 
            .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r [4]), .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r [3]), 
<<<<<<< HEAD
            .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r [2]), .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r [1]), 
            .rx_buf_byte({rx_buf_byte}), .n5734(n5734), .\fifo_temp_output[1] (fifo_temp_output[1]), 
            .n10640(n10640), .VCC_net(VCC_net), .n5738(n5738), .\fifo_temp_output[2] (fifo_temp_output[2]), 
            .n5633(n5633), .rd_fifo_en_prev_r(rd_fifo_en_prev_r), .fifo_read_cmd(fifo_read_cmd), 
            .is_fifo_empty_flag(is_fifo_empty_flag), .empty_o_N_1333(empty_o_N_1333), 
            .n11046(n11046), .n5741(n5741), .\fifo_temp_output[3] (fifo_temp_output[3]), 
            .n5745(n5745), .\fifo_temp_output[4] (fifo_temp_output[4]), 
            .n5748(n5748), .\fifo_temp_output[5] (fifo_temp_output[5]), 
            .n5812(n5812), .\fifo_temp_output[0] (fifo_temp_output[0]), 
            .n5755(n5755), .\fifo_temp_output[6] (fifo_temp_output[6]), 
            .n5761(n5761), .\fifo_temp_output[7] (fifo_temp_output[7]), 
            .n5769(n5769), .n5610(n5610), .n5614(n5614), .\rd_addr_p1_w[2] (rd_addr_p1_w_adj_1495[2]), 
            .n11863(n11863)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(1024[16] 1040[2])
    SB_LUT4 i4164_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5623));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4164_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4362_3_lut (.I0(n5527), .I1(r_Bit_Index[0]), .I2(n5214), 
            .I3(GND_net), .O(n5821));   // src/uart_rx.v(49[10] 144[8])
    defparam i4362_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i4166_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5625));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4166_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4167_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5626));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4167_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut_adj_137 (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(wr_addr_r_adj_1490[0]), .I3(rd_addr_r_adj_1493[0]), .O(n4));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_2_lut_4_lut_adj_137.LUT_INIT = 16'h0220;
    \uart_tx(CLKS_PER_BIT=20)  pc_tx (.r_SM_Main({r_SM_Main_adj_1435}), .\r_SM_Main_2__N_1025[1] (r_SM_Main_2__N_1025[1]), 
            .UART_TX_c(UART_TX_c), .SLM_CLK_c(SLM_CLK_c), .n11691(n11691), 
            .r_Bit_Index({Open_0, Open_1, r_Bit_Index_adj_1437[0]}), .GND_net(GND_net), 
            .n5716(n5716), .r_Tx_Data({r_Tx_Data}), .n5715(n5715), .n5714(n5714), 
            .n5713(n5713), .\r_SM_Main_2__N_1028[0] (r_SM_Main_2__N_1028[0]), 
            .n11079(n11079), .n5712(n5712), .n5711(n5711), .n5710(n5710), 
            .VCC_net(VCC_net), .n5212(n5212), .n5525(n5525), .n5817(n5817), 
            .n5618(n5618), .n5617(n5617), .tx_uart_active_flag(tx_uart_active_flag), 
            .n4715(n4715)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(859[42] 868[3])
    SB_LUT4 i1_4_lut_adj_138 (.I0(rd_addr_r_adj_1493[1]), .I1(rd_addr_r_adj_1493[0]), 
            .I2(wr_addr_r_adj_1490[1]), .I3(wr_addr_r_adj_1490[0]), .O(n32));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_adj_138.LUT_INIT = 16'h8421;
    SB_LUT4 i4240_3_lut (.I0(rx_buf_byte[1]), .I1(rx_shift_reg[1]), .I2(n5120), 
            .I3(GND_net), .O(n5699));   // src/spi.v(76[8] 221[4])
    defparam i4240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4241_3_lut (.I0(rx_shift_reg[7]), .I1(rx_shift_reg[6]), .I2(n5113), 
            .I3(GND_net), .O(n5700));   // src/spi.v(76[8] 221[4])
    defparam i4241_3_lut.LUT_INIT = 16'hcaca;
    fifo_dc_32_lut_gen2 fifo_dc_32_lut_gen_inst (.n30(n30), .n31(n31), .n5731(n5731), 
            .\REG.mem_28_0 (\REG.mem_28_0 ), .FIFO_CLK_c(FIFO_CLK_c), .GND_net(GND_net), 
            .n5726(n5726), .\REG.mem_27_0 (\REG.mem_27_0 ), .n5725(n5725), 
            .\REG.mem_26_0 (\REG.mem_26_0 ), .rd_fifo_en_w(rd_fifo_en_w), 
            .DEBUG_5_c_0(DEBUG_5_c_0), .SLM_CLK_c(SLM_CLK_c), .DEBUG_1_c(DEBUG_1_c), 
            .reset_per_frame(reset_per_frame), .n5723(n5723), .\REG.mem_25_0 (\REG.mem_25_0 ), 
            .\REG.mem_16_0 (\REG.mem_16_0 ), .\REG.mem_17_0 (\REG.mem_17_0 ), 
            .\rd_addr_r[0] (rd_addr_r[0]), .\REG.mem_18_0 (\REG.mem_18_0 ), 
            .\REG.mem_19_0 (\REG.mem_19_0 ), .n5721(n5721), .\REG.mem_24_0 (\REG.mem_24_0 ), 
            .\rd_grey_sync_r[0] (rd_grey_sync_r[0]), .\wr_addr_r[4] (wr_addr_r[4]), 
            .DEBUG_9_c(DEBUG_9_c), .wr_grey_sync_r({wr_grey_sync_r}), .n5719(n5719), 
            .\REG.mem_23_0 (\REG.mem_23_0 ), .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .DEBUG_6_c(DEBUG_6_c), .VCC_net(VCC_net), .n5718(n5718), .\REG.mem_22_0 (\REG.mem_22_0 ), 
            .n5717(n5717), .\REG.mem_21_0 (\REG.mem_21_0 ), .dc32_fifo_full(dc32_fifo_full), 
            .\REG.mem_20_0 (\REG.mem_20_0 ), .\rd_addr_nxt_c_5__N_572[2] (rd_addr_nxt_c_5__N_572[2]), 
            .n5708(n5708), .n5707(n5707), .\REG.mem_14_0 (\REG.mem_14_0 ), 
            .\REG.mem_15_0 (\REG.mem_15_0 ), .\REG.mem_13_0 (\REG.mem_13_0 ), 
            .\REG.mem_12_0 (\REG.mem_12_0 ), .n5691(n5691), .rp_sync1_r({rp_sync1_r}), 
            .n5690(n5690), .n5689(n5689), .n5688(n5688), .n5687(n5687), 
            .n5686(n5686), .n5685(n5685), .n5684(n5684), .n5683(n5683), 
            .n5682(n5682), .n5681(n5681), .n5679(n5679), .n7(n7), .n6(n6), 
            .\REG.mem_2_0 (\REG.mem_2_0 ), .\REG.mem_3_0 (\REG.mem_3_0 ), 
            .\REG.mem_1_0 (\REG.mem_1_0 ), .\REG.mem_0_0 (\REG.mem_0_0 ), 
            .n5677(n5677), .\rd_addr_r[5] (rd_addr_r[5]), .n5675(n5675), 
            .wp_sync1_r({wp_sync1_r}), .n5674(n5674), .n5673(n5673), .n5672(n5672), 
            .n5671(n5671), .\rd_grey_sync_r[4] (rd_grey_sync_r[4]), .\rd_grey_sync_r[3] (rd_grey_sync_r[3]), 
            .\rd_grey_sync_r[2] (rd_grey_sync_r[2]), .\rd_grey_sync_r[1] (rd_grey_sync_r[1]), 
            .n5670(n5670), .n5669(n5669), .n5668(n5668), .n5667(n5667), 
            .n5666(n5666), .n59(n59), .n47(n47), .n5664(n5664), .n5663(n5663), 
            .n5662(n5662), .n5661(n5661), .\wr_addr_nxt_c[0] (wr_addr_nxt_c[0]), 
            .\wr_addr_nxt_c[1] (wr_addr_nxt_c[1]), .n5659(n5659), .\rd_addr_p1_w[0] (rd_addr_p1_w[0]), 
            .n5657(n5657), .n5655(n5655), .\REG.mem_6_0 (\REG.mem_6_0 ), 
            .\REG.mem_7_0 (\REG.mem_7_0 ), .dc32_fifo_read_enable(dc32_fifo_read_enable), 
            .n5645(n5645), .\REG.mem_11_0 (\REG.mem_11_0 ), .\REG.mem_30_0 (\REG.mem_30_0 ), 
            .\REG.mem_31_0 (\REG.mem_31_0 ), .\REG.mem_29_0 (\REG.mem_29_0 ), 
            .\REG.mem_5_0 (\REG.mem_5_0 ), .\REG.mem_4_0 (\REG.mem_4_0 ), 
            .n5642(n5642), .\REG.mem_10_0 (\REG.mem_10_0 ), .n5641(n5641), 
            .\REG.mem_9_0 (\REG.mem_9_0 ), .n5640(n5640), .\REG.mem_8_0 (\REG.mem_8_0 ), 
            .\wr_addr_nxt_c[2] (wr_addr_nxt_c[2]), .\wr_addr_nxt_c[3] (wr_addr_nxt_c[3]), 
            .\wr_addr_nxt_c[4] (wr_addr_nxt_c[4]), .n25(n25_adj_1405), .\wr_grey_w[5] (wr_grey_w[5]), 
            .n5639(n5639), .dc32_fifo_write_enable(dc32_fifo_write_enable), 
            .n5638(n5638), .n5637(n5637), .n5635(n5635), .n5634(n5634), 
            .n26(n26), .n5631(n5631), .n5626(n5626), .n5625(n5625), 
            .n5624(n5624), .n5623(n5623), .n5622(n5622), .n5615(n5615), 
            .n5611(n5611), .\rd_addr_nxt_c_5__N_572[4] (rd_addr_nxt_c_5__N_572[4]), 
            .n5766(n5766), .n5607(n5607), .n24(n24_adj_1404), .n5762(n5762), 
            .n22(n22), .n20(n20), .n5751(n5751), .n5750(n5750), .n5749(n5749), 
            .n23(n23_adj_1402), .n21(n21), .n5742(n5742), .n28(n28), 
            .n34(n34), .n35(n35), .n5735(n5735), .n32(n32_adj_1403), 
            .n33(n33), .n29(n29), .n27(n27)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(579[21] 595[2])
=======
            .rd_addr_r({rd_addr_r_adj_121}), .reset_all_w(reset_all_w), 
            .n8(n8), .wr_addr_r({wr_addr_r_adj_118}), .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r [2]), 
            .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r [1]), .GND_net(GND_net), 
            .\rd_addr_p1_w[2] (rd_addr_p1_w_adj_123[2]), .n14025(n14025), 
            .n6127(n6127), .VCC_net(VCC_net), .\fifo_temp_output[1] (fifo_temp_output[1]), 
            .n10430(n10430), .is_tx_fifo_full_flag(is_tx_fifo_full_flag), 
            .n6088(n6088), .\fifo_temp_output[0] (fifo_temp_output[0]), 
            .\wr_addr_p1_w[2] (wr_addr_p1_w_adj_120[2]), .n1(n1), .n10226(n10226), 
            .n5989(n5989), .n5311(n5311), .\fifo_temp_output[4] (fifo_temp_output[4]), 
            .n5314(n5314), .\fifo_temp_output[5] (fifo_temp_output[5]), 
            .rx_buf_byte({rx_buf_byte}), .n5868(n5868), .n4882(n4882), 
            .\fifo_temp_output[2] (fifo_temp_output[2]), .n4887(n4887), 
            .\fifo_temp_output[3] (fifo_temp_output[3]), .n5536(n5536), 
            .\fifo_temp_output[6] (fifo_temp_output[6]), .n5539(n5539), 
            .\fifo_temp_output[7] (fifo_temp_output[7]), .n10786(n10786), 
            .is_fifo_empty_flag(is_fifo_empty_flag), .n4919(n4919), .n4922(n4922), 
            .fifo_write_cmd(fifo_write_cmd), .wr_fifo_en_w(wr_fifo_en_w), 
            .n4878(n4878), .rd_fifo_en_prev_r(rd_fifo_en_prev_r), .fifo_read_cmd(fifo_read_cmd)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(933[16] 949[2])
    SB_LUT4 i3579_3_lut (.I0(\REG.mem_3_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n62), .I3(GND_net), .O(n4962));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3579_3_lut.LUT_INIT = 16'hcaca;
    spi spi0 (.\tx_data_byte[3] (tx_data_byte[3]), .n2086(n2086), .GND_net(GND_net), 
        .\tx_data_byte[4] (tx_data_byte[4]), .SEN_c_1(SEN_c_1), .SLM_CLK_c(SLM_CLK_c), 
        .\tx_data_byte[5] (tx_data_byte[5]), .SOUT_c(SOUT_c), .n4312(n4312), 
        .\rx_shift_reg[0] (rx_shift_reg[0]), .\tx_data_byte[6] (tx_data_byte[6]), 
        .n4319(n4319), .SDAT_c_15(SDAT_c_15), .\tx_data_byte[7] (tx_data_byte[7]), 
        .tx_addr_byte({tx_addr_byte}), .VCC_net(VCC_net), .n10428(n10428), 
        .\tx_shift_reg[0] (tx_shift_reg[0]), .n6060(n6060), .rx_buf_byte({rx_buf_byte}), 
        .n6059(n6059), .n6058(n6058), .n6057(n6057), .n6056(n6056), 
        .n6055(n6055), .n6054(n6054), .spi_rx_byte_ready(spi_rx_byte_ready), 
        .SCK_c_0(SCK_c_0), .spi_start_transfer_r(spi_start_transfer_r), 
        .n4897(n4897), .n4888(n4888), .\rx_shift_reg[1] (rx_shift_reg[1]), 
        .n4883(n4883), .\rx_shift_reg[2] (rx_shift_reg[2]), .n4877(n4877), 
        .\rx_shift_reg[3] (rx_shift_reg[3]), .n4869(n4869), .\rx_shift_reg[4] (rx_shift_reg[4]), 
        .n4838(n4838), .\rx_shift_reg[5] (rx_shift_reg[5]), .multi_byte_spi_trans_flag_r(multi_byte_spi_trans_flag_r), 
        .n4836(n4836), .\rx_shift_reg[6] (rx_shift_reg[6]), .n4834(n4834), 
        .\rx_shift_reg[7] (rx_shift_reg[7]), .\tx_data_byte[2] (tx_data_byte[2]), 
        .\tx_data_byte[1] (tx_data_byte[1]), .n3495(n3495)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(833[5] 857[2])
    SB_LUT4 i3578_3_lut (.I0(\REG.mem_3_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n62), .I3(GND_net), .O(n4961));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3578_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3518_2_lut_4_lut (.I0(reset_per_frame), .I1(rd_addr_r[0]), 
            .I2(rd_addr_p1_w[0]), .I3(rd_fifo_en_w), .O(n4901));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i3518_2_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i3536_4_lut_4_lut (.I0(reset_all_w), .I1(rd_addr_r_adj_121[1]), 
            .I2(rd_addr_r_adj_121[0]), .I3(rd_fifo_en_w_adj_56), .O(n4919));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i3536_4_lut_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i4153_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[6]), 
            .I2(\mem_LUT.data_raw_r [6]), .I3(n4459), .O(n5536));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4153_4_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4156_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[7]), 
            .I2(\mem_LUT.data_raw_r [7]), .I3(n4459), .O(n5539));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4156_4_lut_4_lut.LUT_INIT = 16'h5044;
    \uart_tx(CLKS_PER_BIT=20)  pc_tx (.UART_TX_c(UART_TX_c), .SLM_CLK_c(SLM_CLK_c), 
            .r_SM_Main({r_SM_Main_adj_95}), .GND_net(GND_net), .\r_SM_Main_2__N_841[1] (r_SM_Main_2__N_841[1]), 
            .\r_SM_Main_2__N_844[0] (r_SM_Main_2__N_844[0]), .n3794(n3794), 
            .VCC_net(VCC_net), .n13865(n13865), .n10805(n10805), .n4890(n4890), 
            .r_Tx_Data({r_Tx_Data}), .n4889(n4889), .tx_uart_active_flag(tx_uart_active_flag), 
            .n5192(n5192), .n5191(n5191), .n5190(n5190), .n5189(n5189), 
            .n5187(n5187), .n5171(n5171), .n5170(n5170)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(768[42] 777[3])
    usb3_if usb3_if_inst (.reset_per_frame(reset_per_frame), .reset_per_frame_latched(reset_per_frame_latched), 
            .SLM_CLK_c(SLM_CLK_c), .DEBUG_3_c(DEBUG_3_c), .DEBUG_2_c(DEBUG_2_c), 
            .FIFO_CLK_c(FIFO_CLK_c), .\dc32_fifo_data_in[0] (dc32_fifo_data_in[0]), 
            .DEBUG_5_c(DEBUG_5_c), .buffer_switch_done(buffer_switch_done), 
            .buffer_switch_done_latched(buffer_switch_done_latched), .VCC_net(VCC_net), 
            .FT_OE_c(FT_OE_c), .n571(n571), .GND_net(GND_net), .n575(n575), 
            .write_to_dc32_fifo_latched_N_425(write_to_dc32_fifo_latched_N_425), 
            .n2352(n2352), .n4911(n4911), .n4910(n4910), .n4907(n4907), 
            .FIFO_D15_c_15(FIFO_D15_c_15), .FIFO_D14_c_14(FIFO_D14_c_14), 
            .FIFO_D13_c_13(FIFO_D13_c_13), .FIFO_D12_c_12(FIFO_D12_c_12), 
            .FIFO_D11_c_11(FIFO_D11_c_11), .FIFO_D10_c_10(FIFO_D10_c_10), 
            .FIFO_D9_c_9(FIFO_D9_c_9), .FIFO_D8_c_8(FIFO_D8_c_8), .FIFO_D7_c_7(FIFO_D7_c_7), 
            .FIFO_D6_c_6(FIFO_D6_c_6), .FIFO_D5_c_5(FIFO_D5_c_5), .FIFO_D4_c_4(FIFO_D4_c_4), 
            .FIFO_D3_c_3(FIFO_D3_c_3), .FIFO_D2_c_2(FIFO_D2_c_2), .FIFO_D1_c_1(FIFO_D1_c_1), 
            .dc32_fifo_almost_full(dc32_fifo_almost_full), .\dc32_fifo_data_in[15] (dc32_fifo_data_in[15]), 
            .\dc32_fifo_data_in[14] (dc32_fifo_data_in[14]), .\dc32_fifo_data_in[13] (dc32_fifo_data_in[13]), 
            .\dc32_fifo_data_in[12] (dc32_fifo_data_in[12]), .\dc32_fifo_data_in[11] (dc32_fifo_data_in[11]), 
            .\dc32_fifo_data_in[10] (dc32_fifo_data_in[10]), .\dc32_fifo_data_in[9] (dc32_fifo_data_in[9]), 
            .\dc32_fifo_data_in[8] (dc32_fifo_data_in[8]), .\dc32_fifo_data_in[7] (dc32_fifo_data_in[7]), 
            .\dc32_fifo_data_in[6] (dc32_fifo_data_in[6]), .\dc32_fifo_data_in[5] (dc32_fifo_data_in[5]), 
            .\dc32_fifo_data_in[4] (dc32_fifo_data_in[4]), .\dc32_fifo_data_in[3] (dc32_fifo_data_in[3]), 
            .\dc32_fifo_data_in[2] (dc32_fifo_data_in[2]), .\dc32_fifo_data_in[1] (dc32_fifo_data_in[1]), 
            .DEBUG_1_c_c(DEBUG_1_c_c), .FT_OE_N_420(FT_OE_N_420)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(513[9] 530[3])
=======
    SB_IO SDAT_pad (.PACKAGE_PIN(SDAT), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SDAT_c_15)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SDAT_pad.PIN_TYPE = 6'b011001;
    defparam SDAT_pad.PULLUP = 1'b0;
    defparam SDAT_pad.NEG_TRIGGER = 1'b0;
    defparam SDAT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UPDATE_pad (.PACKAGE_PIN(UPDATE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(UPDATE_c_3));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UPDATE_pad.PIN_TYPE = 6'b011001;
    defparam UPDATE_pad.PULLUP = 1'b0;
    defparam UPDATE_pad.NEG_TRIGGER = 1'b0;
    defparam UPDATE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO RESET_pad (.PACKAGE_PIN(RESET), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(RESET_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RESET_pad.PIN_TYPE = 6'b011001;
    defparam RESET_pad.PULLUP = 1'b0;
    defparam RESET_pad.NEG_TRIGGER = 1'b0;
    defparam RESET_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SLM_CLK_pad (.PACKAGE_PIN(SLM_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SLM_CLK_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SLM_CLK_pad.PIN_TYPE = 6'b011001;
    defparam SLM_CLK_pad.PULLUP = 1'b0;
    defparam SLM_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam SLM_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INVERT_pad (.PACKAGE_PIN(INVERT), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INVERT_c_4)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INVERT_pad.PIN_TYPE = 6'b011001;
    defparam INVERT_pad.PULLUP = 1'b0;
    defparam INVERT_pad.NEG_TRIGGER = 1'b0;
    defparam INVERT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SYNC_pad (.PACKAGE_PIN(SYNC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SYNC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SYNC_pad.PIN_TYPE = 6'b011001;
    defparam SYNC_pad.PULLUP = 1'b0;
    defparam SYNC_pad.NEG_TRIGGER = 1'b0;
    defparam SYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO VALID_pad (.PACKAGE_PIN(VALID), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam VALID_pad.PIN_TYPE = 6'b011001;
    defparam VALID_pad.PULLUP = 1'b0;
    defparam VALID_pad.NEG_TRIGGER = 1'b0;
    defparam VALID_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA31_pad (.PACKAGE_PIN(DATA31), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA31_c_31));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA31_pad.PIN_TYPE = 6'b011001;
    defparam DATA31_pad.PULLUP = 1'b0;
    defparam DATA31_pad.NEG_TRIGGER = 1'b0;
    defparam DATA31_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA0_pad (.PACKAGE_PIN(DATA0), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_8_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA0_pad.PIN_TYPE = 6'b011001;
    defparam DATA0_pad.PULLUP = 1'b0;
    defparam DATA0_pad.NEG_TRIGGER = 1'b0;
    defparam DATA0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA30_pad (.PACKAGE_PIN(DATA30), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA30_c_30));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA30_pad.PIN_TYPE = 6'b011001;
    defparam DATA30_pad.PULLUP = 1'b0;
    defparam DATA30_pad.NEG_TRIGGER = 1'b0;
    defparam DATA30_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA29_pad (.PACKAGE_PIN(DATA29), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA29_c_29));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA29_pad.PIN_TYPE = 6'b011001;
    defparam DATA29_pad.PULLUP = 1'b0;
    defparam DATA29_pad.NEG_TRIGGER = 1'b0;
    defparam DATA29_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA1_pad (.PACKAGE_PIN(DATA1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA1_c_1));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA1_pad.PIN_TYPE = 6'b011001;
    defparam DATA1_pad.PULLUP = 1'b0;
    defparam DATA1_pad.NEG_TRIGGER = 1'b0;
    defparam DATA1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA28_pad (.PACKAGE_PIN(DATA28), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA28_c_28));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA28_pad.PIN_TYPE = 6'b011001;
    defparam DATA28_pad.PULLUP = 1'b0;
    defparam DATA28_pad.NEG_TRIGGER = 1'b0;
    defparam DATA28_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA27_pad (.PACKAGE_PIN(DATA27), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA27_c_27));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA27_pad.PIN_TYPE = 6'b011001;
    defparam DATA27_pad.PULLUP = 1'b0;
    defparam DATA27_pad.NEG_TRIGGER = 1'b0;
    defparam DATA27_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA2_pad (.PACKAGE_PIN(DATA2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA2_c_2));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA2_pad.PIN_TYPE = 6'b011001;
    defparam DATA2_pad.PULLUP = 1'b0;
    defparam DATA2_pad.NEG_TRIGGER = 1'b0;
    defparam DATA2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA26_pad (.PACKAGE_PIN(DATA26), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA26_c_26));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA26_pad.PIN_TYPE = 6'b011001;
    defparam DATA26_pad.PULLUP = 1'b0;
    defparam DATA26_pad.NEG_TRIGGER = 1'b0;
    defparam DATA26_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA25_pad (.PACKAGE_PIN(DATA25), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA25_c_25));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA25_pad.PIN_TYPE = 6'b011001;
    defparam DATA25_pad.PULLUP = 1'b0;
    defparam DATA25_pad.NEG_TRIGGER = 1'b0;
    defparam DATA25_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA3_pad (.PACKAGE_PIN(DATA3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA3_c_3));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA3_pad.PIN_TYPE = 6'b011001;
    defparam DATA3_pad.PULLUP = 1'b0;
    defparam DATA3_pad.NEG_TRIGGER = 1'b0;
    defparam DATA3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA24_pad (.PACKAGE_PIN(DATA24), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA24_c_24));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA24_pad.PIN_TYPE = 6'b011001;
    defparam DATA24_pad.PULLUP = 1'b0;
    defparam DATA24_pad.NEG_TRIGGER = 1'b0;
    defparam DATA24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA23_pad (.PACKAGE_PIN(DATA23), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA23_c_23));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA23_pad.PIN_TYPE = 6'b011001;
    defparam DATA23_pad.PULLUP = 1'b0;
    defparam DATA23_pad.NEG_TRIGGER = 1'b0;
    defparam DATA23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA4_pad (.PACKAGE_PIN(DATA4), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA4_c_4));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA4_pad.PIN_TYPE = 6'b011001;
    defparam DATA4_pad.PULLUP = 1'b0;
    defparam DATA4_pad.NEG_TRIGGER = 1'b0;
    defparam DATA4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA22_pad (.PACKAGE_PIN(DATA22), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA22_c_22));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA22_pad.PIN_TYPE = 6'b011001;
    defparam DATA22_pad.PULLUP = 1'b0;
    defparam DATA22_pad.NEG_TRIGGER = 1'b0;
    defparam DATA22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA21_pad (.PACKAGE_PIN(DATA21), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA21_c_21));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA21_pad.PIN_TYPE = 6'b011001;
    defparam DATA21_pad.PULLUP = 1'b0;
    defparam DATA21_pad.NEG_TRIGGER = 1'b0;
    defparam DATA21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA5_pad (.PACKAGE_PIN(DATA5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA5_c_5));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA5_pad.PIN_TYPE = 6'b011001;
    defparam DATA5_pad.PULLUP = 1'b0;
    defparam DATA5_pad.NEG_TRIGGER = 1'b0;
    defparam DATA5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA20_pad (.PACKAGE_PIN(DATA20), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA20_c_20));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA20_pad.PIN_TYPE = 6'b011001;
    defparam DATA20_pad.PULLUP = 1'b0;
    defparam DATA20_pad.NEG_TRIGGER = 1'b0;
    defparam DATA20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA19_pad (.PACKAGE_PIN(DATA19), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA19_c_19));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA19_pad.PIN_TYPE = 6'b011001;
    defparam DATA19_pad.PULLUP = 1'b0;
    defparam DATA19_pad.NEG_TRIGGER = 1'b0;
    defparam DATA19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA6_pad (.PACKAGE_PIN(DATA6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA6_c_6));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA6_pad.PIN_TYPE = 6'b011001;
    defparam DATA6_pad.PULLUP = 1'b0;
    defparam DATA6_pad.NEG_TRIGGER = 1'b0;
    defparam DATA6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA18_pad (.PACKAGE_PIN(DATA18), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA18_c_18));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA18_pad.PIN_TYPE = 6'b011001;
    defparam DATA18_pad.PULLUP = 1'b0;
    defparam DATA18_pad.NEG_TRIGGER = 1'b0;
    defparam DATA18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA17_pad (.PACKAGE_PIN(DATA17), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA17_c_17));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA17_pad.PIN_TYPE = 6'b011001;
    defparam DATA17_pad.PULLUP = 1'b0;
    defparam DATA17_pad.NEG_TRIGGER = 1'b0;
    defparam DATA17_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA7_pad (.PACKAGE_PIN(DATA7), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA7_c_7));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA7_pad.PIN_TYPE = 6'b011001;
    defparam DATA7_pad.PULLUP = 1'b0;
    defparam DATA7_pad.NEG_TRIGGER = 1'b0;
    defparam DATA7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA16_pad (.PACKAGE_PIN(DATA16), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA16_c_16));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA16_pad.PIN_TYPE = 6'b011001;
    defparam DATA16_pad.PULLUP = 1'b0;
    defparam DATA16_pad.NEG_TRIGGER = 1'b0;
    defparam DATA16_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA15_pad (.PACKAGE_PIN(DATA15), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA15_c_15));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA15_pad.PIN_TYPE = 6'b011001;
    defparam DATA15_pad.PULLUP = 1'b0;
    defparam DATA15_pad.NEG_TRIGGER = 1'b0;
    defparam DATA15_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA8_pad (.PACKAGE_PIN(DATA8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA8_c_8));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA8_pad.PIN_TYPE = 6'b011001;
    defparam DATA8_pad.PULLUP = 1'b0;
    defparam DATA8_pad.NEG_TRIGGER = 1'b0;
    defparam DATA8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA14_pad (.PACKAGE_PIN(DATA14), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA14_c_14));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA14_pad.PIN_TYPE = 6'b011001;
    defparam DATA14_pad.PULLUP = 1'b0;
    defparam DATA14_pad.NEG_TRIGGER = 1'b0;
    defparam DATA14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA13_pad (.PACKAGE_PIN(DATA13), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA13_c_13));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA13_pad.PIN_TYPE = 6'b011001;
    defparam DATA13_pad.PULLUP = 1'b0;
    defparam DATA13_pad.NEG_TRIGGER = 1'b0;
    defparam DATA13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA12_pad (.PACKAGE_PIN(DATA12), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA12_c_12));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA12_pad.PIN_TYPE = 6'b011001;
    defparam DATA12_pad.PULLUP = 1'b0;
    defparam DATA12_pad.NEG_TRIGGER = 1'b0;
    defparam DATA12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA11_pad (.PACKAGE_PIN(DATA11), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA11_c_11));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA11_pad.PIN_TYPE = 6'b011001;
    defparam DATA11_pad.PULLUP = 1'b0;
    defparam DATA11_pad.NEG_TRIGGER = 1'b0;
    defparam DATA11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA9_pad (.PACKAGE_PIN(DATA9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA9_c_9));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA9_pad.PIN_TYPE = 6'b011001;
    defparam DATA9_pad.PULLUP = 1'b0;
    defparam DATA9_pad.NEG_TRIGGER = 1'b0;
    defparam DATA9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA10_pad (.PACKAGE_PIN(DATA10), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA10_c_10));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA10_pad.PIN_TYPE = 6'b011001;
    defparam DATA10_pad.PULLUP = 1'b0;
    defparam DATA10_pad.NEG_TRIGGER = 1'b0;
    defparam DATA10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_OE_pad (.PACKAGE_PIN(FT_OE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(FT_OE_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_OE_pad.PIN_TYPE = 6'b011001;
    defparam FT_OE_pad.PULLUP = 1'b0;
    defparam FT_OE_pad.NEG_TRIGGER = 1'b0;
    defparam FT_OE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_RD_pad (.PACKAGE_PIN(FT_RD), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(FT_RD_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_RD_pad.PIN_TYPE = 6'b011001;
    defparam FT_RD_pad.PULLUP = 1'b0;
    defparam FT_RD_pad.NEG_TRIGGER = 1'b0;
    defparam FT_RD_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_WR_pad (.PACKAGE_PIN(FT_WR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_WR_pad.PIN_TYPE = 6'b011001;
    defparam FT_WR_pad.PULLUP = 1'b0;
    defparam FT_WR_pad.NEG_TRIGGER = 1'b0;
    defparam FT_WR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_SIWU_pad (.PACKAGE_PIN(FT_SIWU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_SIWU_pad.PIN_TYPE = 6'b011001;
    defparam FT_SIWU_pad.PULLUP = 1'b0;
    defparam FT_SIWU_pad.NEG_TRIGGER = 1'b0;
    defparam FT_SIWU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_0_pad (.PACKAGE_PIN(DEBUG_0), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_0_c_24));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_0_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_0_pad.PULLUP = 1'b0;
    defparam DEBUG_0_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_1_pad (.PACKAGE_PIN(DEBUG_1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_1_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_1_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_1_pad.PULLUP = 1'b0;
    defparam DEBUG_1_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_2_pad (.PACKAGE_PIN(DEBUG_2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_2_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_2_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_2_pad.PULLUP = 1'b0;
    defparam DEBUG_2_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_3_pad (.PACKAGE_PIN(DEBUG_3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_3_c_0_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_3_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_3_pad.PULLUP = 1'b0;
    defparam DEBUG_3_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_5_pad (.PACKAGE_PIN(DEBUG_5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_5_c_0));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_5_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_5_pad.PULLUP = 1'b0;
    defparam DEBUG_5_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_6_pad (.PACKAGE_PIN(DEBUG_6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_6_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_6_pad.PULLUP = 1'b0;
    defparam DEBUG_6_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_8_pad (.PACKAGE_PIN(DEBUG_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_8_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_8_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_8_pad.PULLUP = 1'b0;
    defparam DEBUG_8_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_9_pad (.PACKAGE_PIN(DEBUG_9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_9_c_0));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_9_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_9_pad.PULLUP = 1'b0;
    defparam DEBUG_9_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CLK_pad (.PACKAGE_PIN(ICE_CLK), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CLK_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CLK_pad.PULLUP = 1'b0;
    defparam ICE_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CDONE_pad (.PACKAGE_PIN(ICE_CDONE), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CDONE_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CDONE_pad.PULLUP = 1'b0;
    defparam ICE_CDONE_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CDONE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CREST_pad (.PACKAGE_PIN(ICE_CREST), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CREST_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CREST_pad.PULLUP = 1'b0;
    defparam ICE_CREST_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CREST_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY led_counter_1434_1494_add_4_24 (.CI(n12175), .I0(GND_net), 
            .I1(n3), .CO(n12176));
    SB_IO ICE_SYSCLK_pad (.PACKAGE_PIN(ICE_SYSCLK), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ICE_SYSCLK_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_SYSCLK_pad.PIN_TYPE = 6'b000001;
    defparam ICE_SYSCLK_pad.PULLUP = 1'b0;
    defparam ICE_SYSCLK_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_SYSCLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UART_RX_pad (.PACKAGE_PIN(UART_RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(UART_RX_c)) /* synthesis IO_FF_IN=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UART_RX_pad.PIN_TYPE = 6'b000001;
    defparam UART_RX_pad.PULLUP = 1'b0;
    defparam UART_RX_pad.NEG_TRIGGER = 1'b0;
    defparam UART_RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SOUT_pad (.PACKAGE_PIN(SOUT), .OUTPUT_ENABLE(VCC_net), .D_IN_0(SOUT_c)) /* synthesis IO_FF_IN=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SOUT_pad.PIN_TYPE = 6'b000001;
    defparam SOUT_pad.PULLUP = 1'b0;
    defparam SOUT_pad.NEG_TRIGGER = 1'b0;
    defparam SOUT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FR_RXF_pad (.PACKAGE_PIN(FR_RXF), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FR_RXF_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FR_RXF_pad.PIN_TYPE = 6'b000001;
    defparam FR_RXF_pad.PULLUP = 1'b0;
    defparam FR_RXF_pad.NEG_TRIGGER = 1'b0;
    defparam FR_RXF_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D31_pad (.PACKAGE_PIN(FIFO_D31), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D31_c_31));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D31_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D31_pad.PULLUP = 1'b0;
    defparam FIFO_D31_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D31_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D30_pad (.PACKAGE_PIN(FIFO_D30), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D30_c_30));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D30_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D30_pad.PULLUP = 1'b0;
    defparam FIFO_D30_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D30_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D29_pad (.PACKAGE_PIN(FIFO_D29), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D29_c_29));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D29_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D29_pad.PULLUP = 1'b0;
    defparam FIFO_D29_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D29_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D28_pad (.PACKAGE_PIN(FIFO_D28), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D28_c_28));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D28_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D28_pad.PULLUP = 1'b0;
    defparam FIFO_D28_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D28_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D27_pad (.PACKAGE_PIN(FIFO_D27), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D27_c_27));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D27_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D27_pad.PULLUP = 1'b0;
    defparam FIFO_D27_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D27_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO FIFO_CLK_pad (.PACKAGE_PIN(FIFO_CLK), .OUTPUT_ENABLE(VCC_net), 
            .GLOBAL_BUFFER_OUTPUT(FIFO_CLK_c));   // src/top.v(84[12:20])
    defparam FIFO_CLK_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_CLK_pad.PULLUP = 1'b0;
    defparam FIFO_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D26_pad (.PACKAGE_PIN(FIFO_D26), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D26_c_26));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D26_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D26_pad.PULLUP = 1'b0;
    defparam FIFO_D26_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D26_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D25_pad (.PACKAGE_PIN(FIFO_D25), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D25_c_25));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D25_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D25_pad.PULLUP = 1'b0;
    defparam FIFO_D25_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D25_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D24_pad (.PACKAGE_PIN(FIFO_D24), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D24_c_24));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D24_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D24_pad.PULLUP = 1'b0;
    defparam FIFO_D24_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D23_pad (.PACKAGE_PIN(FIFO_D23), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D23_c_23));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D23_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D23_pad.PULLUP = 1'b0;
    defparam FIFO_D23_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D22_pad (.PACKAGE_PIN(FIFO_D22), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D22_c_22));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D22_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D22_pad.PULLUP = 1'b0;
    defparam FIFO_D22_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D21_pad (.PACKAGE_PIN(FIFO_D21), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D21_c_21));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D21_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D21_pad.PULLUP = 1'b0;
    defparam FIFO_D21_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D20_pad (.PACKAGE_PIN(FIFO_D20), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D20_c_20));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D20_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D20_pad.PULLUP = 1'b0;
    defparam FIFO_D20_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D19_pad (.PACKAGE_PIN(FIFO_D19), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D19_c_19));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D19_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D19_pad.PULLUP = 1'b0;
    defparam FIFO_D19_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D18_pad (.PACKAGE_PIN(FIFO_D18), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D18_c_18));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D18_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D18_pad.PULLUP = 1'b0;
    defparam FIFO_D18_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D17_pad (.PACKAGE_PIN(FIFO_D17), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D17_c_17));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D17_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D17_pad.PULLUP = 1'b0;
    defparam FIFO_D17_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D17_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D16_pad (.PACKAGE_PIN(FIFO_D16), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D16_c_16));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D16_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D16_pad.PULLUP = 1'b0;
    defparam FIFO_D16_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D16_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D15_pad (.PACKAGE_PIN(FIFO_D15), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D15_c_15));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D15_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D15_pad.PULLUP = 1'b0;
    defparam FIFO_D15_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D15_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D14_pad (.PACKAGE_PIN(FIFO_D14), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D14_c_14));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D14_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D14_pad.PULLUP = 1'b0;
    defparam FIFO_D14_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D13_pad (.PACKAGE_PIN(FIFO_D13), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D13_c_13));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D13_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D13_pad.PULLUP = 1'b0;
    defparam FIFO_D13_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D12_pad (.PACKAGE_PIN(FIFO_D12), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D12_c_12));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D12_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D12_pad.PULLUP = 1'b0;
    defparam FIFO_D12_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D11_pad (.PACKAGE_PIN(FIFO_D11), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D11_c_11));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D11_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D11_pad.PULLUP = 1'b0;
    defparam FIFO_D11_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D10_pad (.PACKAGE_PIN(FIFO_D10), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D10_c_10));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D10_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D10_pad.PULLUP = 1'b0;
    defparam FIFO_D10_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D9_pad (.PACKAGE_PIN(FIFO_D9), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D9_c_9));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D9_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D9_pad.PULLUP = 1'b0;
    defparam FIFO_D9_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D8_pad (.PACKAGE_PIN(FIFO_D8), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D8_c_8));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D8_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D8_pad.PULLUP = 1'b0;
    defparam FIFO_D8_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D7_pad (.PACKAGE_PIN(FIFO_D7), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D7_c_7));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D7_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D7_pad.PULLUP = 1'b0;
    defparam FIFO_D7_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D6_pad (.PACKAGE_PIN(FIFO_D6), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D6_c_6));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D6_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D6_pad.PULLUP = 1'b0;
    defparam FIFO_D6_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D5_pad (.PACKAGE_PIN(FIFO_D5), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D5_c_5));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D5_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D5_pad.PULLUP = 1'b0;
    defparam FIFO_D5_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D4_pad (.PACKAGE_PIN(FIFO_D4), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D4_c_4));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D4_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D4_pad.PULLUP = 1'b0;
    defparam FIFO_D4_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D3_pad (.PACKAGE_PIN(FIFO_D3), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D3_c_3));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D3_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D3_pad.PULLUP = 1'b0;
    defparam FIFO_D3_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D2_pad (.PACKAGE_PIN(FIFO_D2), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D2_c_2));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D2_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D2_pad.PULLUP = 1'b0;
    defparam FIFO_D2_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D1_pad (.PACKAGE_PIN(FIFO_D1), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D1_c_1));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D1_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D1_pad.PULLUP = 1'b0;
    defparam FIFO_D1_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_3_c_0_pad (.PACKAGE_PIN(FIFO_D0), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(DEBUG_3_c_0_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_3_c_0_pad.PIN_TYPE = 6'b000001;
    defparam DEBUG_3_c_0_pad.PULLUP = 1'b0;
    defparam DEBUG_3_c_0_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_3_c_0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4910_3_lut (.I0(\REG.mem_24_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n9), .I3(GND_net), .O(n6384));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4910_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR multi_byte_spi_trans_flag_r_86 (.Q(multi_byte_spi_trans_flag_r), 
            .C(SLM_CLK_c), .D(multi_byte_spi_trans_flag_r_N_72), .R(n5384));   // src/top.v(1165[8] 1232[4])
    SB_LUT4 i4911_3_lut (.I0(\REG.mem_24_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n9), .I3(GND_net), .O(n6385));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1434_1494_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4), .I3(n12174), .O(n109)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_23 (.CI(n12174), .I0(GND_net), 
            .I1(n4), .CO(n12175));
    SB_LUT4 led_counter_1434_1494_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5), .I3(n12173), .O(n110)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_22 (.CI(n12173), .I0(GND_net), 
            .I1(n5), .CO(n12174));
    SB_LUT4 led_counter_1434_1494_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_1433), .I3(n12172), .O(n111)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_21 (.CI(n12172), .I0(GND_net), 
            .I1(n6_adj_1433), .CO(n12173));
    SB_LUT4 led_counter_1434_1494_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_1432), .I3(n12171), .O(n112)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_20 (.CI(n12171), .I0(GND_net), 
            .I1(n7_adj_1432), .CO(n12172));
    SB_LUT4 led_counter_1434_1494_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_1431), .I3(n12170), .O(n113)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_19 (.CI(n12170), .I0(GND_net), 
            .I1(n8_adj_1431), .CO(n12171));
    SB_LUT4 i4912_3_lut (.I0(\REG.mem_24_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n9), .I3(GND_net), .O(n6386));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4913_3_lut (.I0(\REG.mem_24_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n9), .I3(GND_net), .O(n6387));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4914_3_lut (.I0(\REG.mem_24_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n9), .I3(GND_net), .O(n6388));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4915_3_lut (.I0(\REG.mem_24_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n9), .I3(GND_net), .O(n6389));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1434_1494_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_1430), .I3(n12169), .O(n114)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4916_3_lut (.I0(\REG.mem_24_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n9), .I3(GND_net), .O(n6390));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4917_3_lut (.I0(\REG.mem_24_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n9), .I3(GND_net), .O(n6391));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4917_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1434_1494_add_4_18 (.CI(n12169), .I0(GND_net), 
            .I1(n9_adj_1430), .CO(n12170));
    SB_LUT4 led_counter_1434_1494_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_1429), .I3(n12168), .O(n115)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_17 (.CI(n12168), .I0(GND_net), 
            .I1(n10_adj_1429), .CO(n12169));
    SB_LUT4 led_counter_1434_1494_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_1428), .I3(n12167), .O(n116)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_16 (.CI(n12167), .I0(GND_net), 
            .I1(n11_adj_1428), .CO(n12168));
    SB_LUT4 led_counter_1434_1494_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_1427), .I3(n12166), .O(n117)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_15 (.CI(n12166), .I0(GND_net), 
            .I1(n12_adj_1427), .CO(n12167));
    SB_LUT4 led_counter_1434_1494_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_1426), .I3(n12165), .O(n118)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4918_3_lut (.I0(\REG.mem_24_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n9), .I3(GND_net), .O(n6392));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4919_3_lut (.I0(\REG.mem_24_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n9), .I3(GND_net), .O(n6393));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4920_3_lut (.I0(\REG.mem_24_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n9), .I3(GND_net), .O(n6394));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4921_3_lut (.I0(\REG.mem_24_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n9), .I3(GND_net), .O(n6395));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4922_3_lut (.I0(\REG.mem_24_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n9), .I3(GND_net), .O(n6396));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4923_3_lut (.I0(\REG.mem_24_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n9), .I3(GND_net), .O(n6397));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4924_3_lut (.I0(\REG.mem_25_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6398));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4925_3_lut (.I0(\REG.mem_25_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6399));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4926_3_lut (.I0(\REG.mem_25_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6400));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4927_3_lut (.I0(\REG.mem_25_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6401));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4928_3_lut (.I0(\REG.mem_25_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6402));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4929_3_lut (.I0(\REG.mem_25_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6403));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4930_3_lut (.I0(\REG.mem_25_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6404));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4930_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF fifo_write_cmd_79 (.Q(fifo_write_cmd), .C(SLM_CLK_c), .D(n5635));   // src/top.v(980[8] 989[4])
    SB_LUT4 i4931_3_lut (.I0(\REG.mem_25_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6405));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4932_3_lut (.I0(\REG.mem_25_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6406));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4933_3_lut (.I0(\REG.mem_25_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6407));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4934_3_lut (.I0(\REG.mem_25_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6408));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4935_3_lut (.I0(\REG.mem_25_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6409));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4936_3_lut (.I0(\REG.mem_25_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6410));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4937_3_lut (.I0(\REG.mem_25_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6411));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4938_3_lut (.I0(\REG.mem_25_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6412));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4939_3_lut (.I0(\REG.mem_25_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6413));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4940_3_lut (.I0(\REG.mem_25_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6414));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4940_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1434_1494_add_4_14 (.CI(n12165), .I0(GND_net), 
            .I1(n13_adj_1426), .CO(n12166));
    SB_LUT4 led_counter_1434_1494_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14), .I3(n12164), .O(n119)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_13 (.CI(n12164), .I0(GND_net), 
            .I1(n14), .CO(n12165));
    SB_LUT4 led_counter_1434_1494_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_1425), .I3(n12163), .O(n120)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_12 (.CI(n12163), .I0(GND_net), 
            .I1(n15_adj_1425), .CO(n12164));
    SB_LUT4 led_counter_1434_1494_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_1424), .I3(n12162), .O(n121)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_11 (.CI(n12162), .I0(GND_net), 
            .I1(n16_adj_1424), .CO(n12163));
    SB_LUT4 led_counter_1434_1494_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17), .I3(n12161), .O(n122)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_10 (.CI(n12161), .I0(GND_net), 
            .I1(n17), .CO(n12162));
    SB_LUT4 led_counter_1434_1494_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18), .I3(n12160), .O(n123)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4941_3_lut (.I0(\REG.mem_25_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6415));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4941_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1434_1494_add_4_9 (.CI(n12160), .I0(GND_net), .I1(n18), 
            .CO(n12161));
    SB_LUT4 led_counter_1434_1494_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19), .I3(n12159), .O(n124)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_8 (.CI(n12159), .I0(GND_net), .I1(n19), 
            .CO(n12160));
    SB_LUT4 led_counter_1434_1494_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20), .I3(n12158), .O(n125)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_7 (.CI(n12158), .I0(GND_net), .I1(n20), 
            .CO(n12159));
    SB_LUT4 led_counter_1434_1494_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21), .I3(n12157), .O(n126)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4668_3_lut (.I0(\REG.mem_17_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n16), .I3(GND_net), .O(n6142));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4669_3_lut (.I0(\REG.mem_17_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n16), .I3(GND_net), .O(n6143));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4670_3_lut (.I0(\REG.mem_17_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n16), .I3(GND_net), .O(n6144));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4671_3_lut (.I0(\REG.mem_17_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n16), .I3(GND_net), .O(n6145));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4672_3_lut (.I0(\REG.mem_17_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n16), .I3(GND_net), .O(n6146));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4673_3_lut (.I0(\REG.mem_17_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n16), .I3(GND_net), .O(n6147));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4942_3_lut (.I0(\REG.mem_25_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6416));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4674_3_lut (.I0(\REG.mem_17_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n16), .I3(GND_net), .O(n6148));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4675_3_lut (.I0(\REG.mem_17_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n16), .I3(GND_net), .O(n6149));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4943_3_lut (.I0(\REG.mem_25_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6417));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4944_3_lut (.I0(\REG.mem_25_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6418));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4945_3_lut (.I0(\REG.mem_25_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6419));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4945_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1434_1494_add_4_6 (.CI(n12157), .I0(GND_net), .I1(n21), 
            .CO(n12158));
    SB_LUT4 led_counter_1434_1494_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_1423), .I3(n12156), .O(n127)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_5 (.CI(n12156), .I0(GND_net), .I1(n22_adj_1423), 
            .CO(n12157));
    SB_LUT4 led_counter_1434_1494_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_1422), .I3(n12155), .O(n128)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1434_1494_add_4_4 (.CI(n12155), .I0(GND_net), .I1(n23_adj_1422), 
            .CO(n12156));
    SB_LUT4 led_counter_1434_1494_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_1421), .I3(n12154), .O(n129)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4946_3_lut (.I0(\REG.mem_25_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6420));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4947_3_lut (.I0(\REG.mem_25_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6421));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4948_3_lut (.I0(\REG.mem_25_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6422));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4949_3_lut (.I0(\REG.mem_25_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6423));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4950_3_lut (.I0(\REG.mem_25_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6424));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4951_3_lut (.I0(\REG.mem_25_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6425));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4952_3_lut (.I0(\REG.mem_25_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6426));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4676_3_lut (.I0(\REG.mem_17_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n16), .I3(GND_net), .O(n6150));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4953_3_lut (.I0(\REG.mem_25_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6427));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4954_3_lut (.I0(\REG.mem_25_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6428));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4677_3_lut (.I0(\REG.mem_17_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n16), .I3(GND_net), .O(n6151));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4678_3_lut (.I0(\REG.mem_17_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n16), .I3(GND_net), .O(n6152));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4679_3_lut (.I0(\REG.mem_17_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n16), .I3(GND_net), .O(n6153));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4680_3_lut (.I0(\REG.mem_17_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n16), .I3(GND_net), .O(n6154));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4681_3_lut (.I0(\REG.mem_17_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n16), .I3(GND_net), .O(n6155));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4682_3_lut (.I0(\REG.mem_17_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n16), .I3(GND_net), .O(n6156));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4682_3_lut.LUT_INIT = 16'hcaca;
    GND i1 (.Y(GND_net));
    SB_LUT4 i4683_3_lut (.I0(\REG.mem_17_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n16), .I3(GND_net), .O(n6157));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4955_3_lut (.I0(\REG.mem_25_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n8_adj_1419), .I3(GND_net), .O(n6429));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4956_3_lut (.I0(\REG.mem_26_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n7), .I3(GND_net), .O(n6430));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4684_3_lut (.I0(\REG.mem_17_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n16), .I3(GND_net), .O(n6158));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4684_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1434_1494_add_4_3 (.CI(n12154), .I0(GND_net), .I1(n24_adj_1421), 
            .CO(n12155));
    SB_LUT4 i4957_3_lut (.I0(\REG.mem_26_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n7), .I3(GND_net), .O(n6431));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4958_3_lut (.I0(\REG.mem_26_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n7), .I3(GND_net), .O(n6432));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4959_3_lut (.I0(\REG.mem_26_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n7), .I3(GND_net), .O(n6433));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4960_3_lut (.I0(\REG.mem_26_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n7), .I3(GND_net), .O(n6434));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4961_3_lut (.I0(\REG.mem_26_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n7), .I3(GND_net), .O(n6435));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4962_3_lut (.I0(\REG.mem_26_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n7), .I3(GND_net), .O(n6436));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4963_3_lut (.I0(\REG.mem_26_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n7), .I3(GND_net), .O(n6437));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4964_3_lut (.I0(\REG.mem_26_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n7), .I3(GND_net), .O(n6438));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4965_3_lut (.I0(\REG.mem_26_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n7), .I3(GND_net), .O(n6439));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4966_3_lut (.I0(\REG.mem_26_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n7), .I3(GND_net), .O(n6440));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4967_3_lut (.I0(\REG.mem_26_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n7), .I3(GND_net), .O(n6441));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4968_3_lut (.I0(\REG.mem_26_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n7), .I3(GND_net), .O(n6442));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4969_3_lut (.I0(\REG.mem_26_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n7), .I3(GND_net), .O(n6443));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4969_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4970_3_lut (.I0(\REG.mem_26_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n7), .I3(GND_net), .O(n6444));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4971_3_lut (.I0(\REG.mem_26_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n7), .I3(GND_net), .O(n6445));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4972_3_lut (.I0(\REG.mem_26_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n7), .I3(GND_net), .O(n6446));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4972_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_addr_byte_r_i0_i0 (.Q(tx_addr_byte[0]), .C(SLM_CLK_c), .D(n5615));   // src/top.v(1165[8] 1232[4])
    SB_LUT4 i4685_3_lut (.I0(\REG.mem_17_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n16), .I3(GND_net), .O(n6159));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4686_3_lut (.I0(\REG.mem_17_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n16), .I3(GND_net), .O(n6160));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4687_3_lut (.I0(\REG.mem_17_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n16), .I3(GND_net), .O(n6161));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4688_3_lut (.I0(\REG.mem_17_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n16), .I3(GND_net), .O(n6162));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4689_3_lut (.I0(\REG.mem_17_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n16), .I3(GND_net), .O(n6163));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4690_3_lut (.I0(\REG.mem_17_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n16), .I3(GND_net), .O(n6164));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4691_3_lut (.I0(\REG.mem_17_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n16), .I3(GND_net), .O(n6165));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4692_3_lut (.I0(\REG.mem_17_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n16), .I3(GND_net), .O(n6166));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4693_3_lut (.I0(\REG.mem_17_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n16), .I3(GND_net), .O(n6167));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3694_4_lut (.I0(n63), .I1(n4688), .I2(n9015), .I3(state[3]), 
            .O(n2075));   // src/timing_controller.v(78[11:16])
    defparam i3694_4_lut.LUT_INIT = 16'h0a88;
    SB_LUT4 i4694_3_lut (.I0(\REG.mem_17_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n16), .I3(GND_net), .O(n6168));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4694_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1434_1494__i1 (.Q(n24_adj_1421), .C(SLM_CLK_c), .D(n129));   // src/top.v(203[20:35])
    SB_LUT4 i4695_3_lut (.I0(\REG.mem_17_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n16), .I3(GND_net), .O(n6169));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4696_3_lut (.I0(\REG.mem_17_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n16), .I3(GND_net), .O(n6170));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4697_3_lut (.I0(\REG.mem_17_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n16), .I3(GND_net), .O(n6171));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4698_3_lut (.I0(\REG.mem_17_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n16), .I3(GND_net), .O(n6172));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4125_4_lut_4_lut (.I0(wr_fifo_en_w_adj_1416), .I1(reset_all_w), 
            .I2(wr_addr_p1_w_adj_1519[2]), .I3(wr_addr_r_adj_1517[2]), .O(n5599));
    defparam i4125_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4133_4_lut_4_lut_4_lut (.I0(wr_fifo_en_w_adj_1416), .I1(reset_all_w), 
            .I2(wr_addr_r_adj_1517[0]), .I3(wr_addr_r_adj_1517[1]), .O(n5607));
    defparam i4133_4_lut_4_lut_4_lut.LUT_INIT = 16'h1320;
    SB_DFF reset_all_r_77 (.Q(reset_all_w), .C(SLM_CLK_c), .D(reset_all_w_N_61));   // src/top.v(246[8] 264[4])
    SB_LUT4 i1_2_lut_adj_123 (.I0(state[3]), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n12906));   // src/timing_controller.v(154[8] 230[4])
    defparam i1_2_lut_adj_123.LUT_INIT = 16'hbbbb;
    SB_LUT4 i5429_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[7]), .I2(r_Bit_Index[0]), 
            .I3(n4787), .O(n6903));   // src/uart_rx.v(49[10] 144[8])
    defparam i5429_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i5430_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[6]), .I2(r_Bit_Index[0]), 
            .I3(n4787), .O(n6904));   // src/uart_rx.v(49[10] 144[8])
    defparam i5430_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i5431_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[5]), .I2(n4_adj_1434), 
            .I3(n4794), .O(n6905));   // src/uart_rx.v(49[10] 144[8])
    defparam i5431_4_lut.LUT_INIT = 16'hccca;
    SB_DFF uart_rx_complete_rising_edge_82 (.Q(uart_rx_complete_rising_edge), 
           .C(SLM_CLK_c), .D(n5592));   // src/top.v(1156[8] 1162[4])
    SB_LUT4 i5432_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[4]), .I2(n4_adj_1434), 
            .I3(n4790), .O(n6906));   // src/uart_rx.v(49[10] 144[8])
    defparam i5432_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i5433_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[3]), .I2(n4_adj_1436), 
            .I3(n4794), .O(n6907));   // src/uart_rx.v(49[10] 144[8])
    defparam i5433_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4699_3_lut (.I0(\REG.mem_17_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n16), .I3(GND_net), .O(n6173));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1434_1494_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_1437), .I3(VCC_net), .O(n130)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1434_1494_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5434_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[2]), .I2(n4_adj_1436), 
            .I3(n4790), .O(n6908));   // src/uart_rx.v(49[10] 144[8])
    defparam i5434_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i5435_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[1]), .I2(n4_adj_1435), 
            .I3(n4794), .O(n6909));   // src/uart_rx.v(49[10] 144[8])
    defparam i5435_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY led_counter_1434_1494_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(n25_adj_1437), .CO(n12154));
    SB_LUT4 i7544_3_lut (.I0(state[1]), .I1(n63), .I2(state[0]), .I3(GND_net), 
            .O(n9013));
    defparam i7544_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i1_3_lut (.I0(state[2]), .I1(state[1]), .I2(state[0]), .I3(GND_net), 
            .O(n4688));   // src/timing_controller.v(78[11:16])
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF led_counter_1434_1494__i2 (.Q(n23_adj_1422), .C(SLM_CLK_c), .D(n128));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i3 (.Q(n22_adj_1423), .C(SLM_CLK_c), .D(n127));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i4 (.Q(n21), .C(SLM_CLK_c), .D(n126));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i5 (.Q(n20), .C(SLM_CLK_c), .D(n125));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i6 (.Q(n19), .C(SLM_CLK_c), .D(n124));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i7 (.Q(n18), .C(SLM_CLK_c), .D(n123));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i8 (.Q(n17), .C(SLM_CLK_c), .D(n122));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i9 (.Q(n16_adj_1424), .C(SLM_CLK_c), .D(n121));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i10 (.Q(n15_adj_1425), .C(SLM_CLK_c), 
           .D(n120));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i11 (.Q(n14), .C(SLM_CLK_c), .D(n119));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i12 (.Q(n13_adj_1426), .C(SLM_CLK_c), 
           .D(n118));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i13 (.Q(n12_adj_1427), .C(SLM_CLK_c), 
           .D(n117));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i14 (.Q(n11_adj_1428), .C(SLM_CLK_c), 
           .D(n116));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i15 (.Q(n10_adj_1429), .C(SLM_CLK_c), 
           .D(n115));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i16 (.Q(n9_adj_1430), .C(SLM_CLK_c), .D(n114));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i17 (.Q(n8_adj_1431), .C(SLM_CLK_c), .D(n113));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i18 (.Q(n7_adj_1432), .C(SLM_CLK_c), .D(n112));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i19 (.Q(n6_adj_1433), .C(SLM_CLK_c), .D(n111));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i20 (.Q(n5), .C(SLM_CLK_c), .D(n110));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i21 (.Q(n4), .C(SLM_CLK_c), .D(n109));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i22 (.Q(n3), .C(SLM_CLK_c), .D(n108));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i23 (.Q(n2), .C(SLM_CLK_c), .D(n107));   // src/top.v(203[20:35])
    SB_DFF led_counter_1434_1494__i24 (.Q(DEBUG_0_c_24), .C(SLM_CLK_c), 
           .D(n106));   // src/top.v(203[20:35])
    SB_DFF reset_clk_counter_i3_1435__i1 (.Q(reset_clk_counter[1]), .C(SLM_CLK_c), 
           .D(n12310));   // src/top.v(259[27:51])
    SB_LUT4 i19_4_lut (.I0(n4688), .I1(n14242), .I2(state[3]), .I3(n63), 
            .O(n12477));   // src/timing_controller.v(154[8] 230[4])
    defparam i19_4_lut.LUT_INIT = 16'hfcac;
    SB_LUT4 i1_2_lut_3_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(reset_clk_counter[1]), .I3(GND_net), .O(n12310));   // src/top.v(259[27:51])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_DFF reset_clk_counter_i3_1435__i2 (.Q(reset_clk_counter[2]), .C(SLM_CLK_c), 
           .D(n12304));   // src/top.v(259[27:51])
    SB_LUT4 i10079_2_lut_3_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(reset_clk_counter[1]), .I3(GND_net), .O(n12040));   // src/top.v(259[27:51])
    defparam i10079_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_DFF reset_clk_counter_i3_1435__i3 (.Q(reset_clk_counter[3]), .C(SLM_CLK_c), 
           .D(n12308));   // src/top.v(259[27:51])
    SB_LUT4 i5454_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6928));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i5454_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1119_4_lut (.I0(n2335), .I1(n9015), .I2(state[3]), .I3(n63), 
            .O(n2180));   // src/timing_controller.v(78[11:16])
    defparam i1119_4_lut.LUT_INIT = 16'h0a3a;
    SB_DFF tx_data_byte_r_i0_i0 (.Q(tx_data_byte[0]), .C(SLM_CLK_c), .D(n5552));   // src/top.v(1165[8] 1232[4])
    SB_LUT4 i5456_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6930));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i5456_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5458_3_lut (.I0(tx_data_byte[7]), .I1(pc_data_rx[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6932));   // src/top.v(1165[8] 1232[4])
    defparam i5458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5459_3_lut (.I0(tx_data_byte[6]), .I1(pc_data_rx[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6933));   // src/top.v(1165[8] 1232[4])
    defparam i5459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5460_3_lut (.I0(tx_data_byte[5]), .I1(pc_data_rx[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6934));   // src/top.v(1165[8] 1232[4])
    defparam i5460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5461_3_lut (.I0(tx_data_byte[4]), .I1(pc_data_rx[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6935));   // src/top.v(1165[8] 1232[4])
    defparam i5461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5462_3_lut (.I0(tx_data_byte[3]), .I1(pc_data_rx[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6936));   // src/top.v(1165[8] 1232[4])
    defparam i5462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5463_3_lut (.I0(tx_data_byte[2]), .I1(pc_data_rx[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6937));   // src/top.v(1165[8] 1232[4])
    defparam i5463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5464_3_lut (.I0(tx_data_byte[1]), .I1(pc_data_rx[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6938));   // src/top.v(1165[8] 1232[4])
    defparam i5464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4191_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[1]), .I2(\mem_LUT.data_raw_r [1]), 
            .I3(n5086), .O(n5665));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4191_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4188_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[2]), .I2(\mem_LUT.data_raw_r [2]), 
            .I3(n5086), .O(n5662));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4188_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i2017_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n3468));   // src/top.v(1165[8] 1232[4])
    defparam i2017_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4185_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[3]), .I2(\mem_LUT.data_raw_r [3]), 
            .I3(n5086), .O(n5659));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4185_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i12300_2_lut (.I0(is_fifo_empty_flag), .I1(tx_uart_active_flag), 
            .I2(GND_net), .I3(GND_net), .O(start_tx_N_64));
    defparam i12300_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i4182_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[4]), .I2(\mem_LUT.data_raw_r [4]), 
            .I3(n5086), .O(n5656));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4182_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i5473_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[0]), .I2(\mem_LUT.data_raw_r [0]), 
            .I3(n5086), .O(n6947));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i5473_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4080_2_lut_4_lut (.I0(reset_per_frame), .I1(wr_addr_r[0]), 
            .I2(wr_addr_p1_w[0]), .I3(wr_fifo_en_w), .O(n5554));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4080_2_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4101_4_lut_4_lut (.I0(tx_uart_active_flag), .I1(r_SM_Main_adj_1467[1]), 
            .I2(r_SM_Main_adj_1467[2]), .I3(n4_adj_1442), .O(n5575));   // src/uart_tx.v(38[10] 141[8])
    defparam i4101_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i1_2_lut_4_lut (.I0(reset_clk_counter[2]), .I1(reset_all_w_N_61), 
            .I2(reset_clk_counter[0]), .I3(reset_clk_counter[1]), .O(n12304));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'haaa6;
    SB_LUT4 i1_2_lut_4_lut_adj_124 (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(wr_addr_r_adj_1517[0]), .I3(rd_addr_r_adj_1520[0]), .O(n4_adj_1441));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_2_lut_4_lut_adj_124.LUT_INIT = 16'h0220;
    SB_LUT4 i4764_3_lut (.I0(\REG.mem_20_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n13), .I3(GND_net), .O(n6238));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4765_3_lut (.I0(\REG.mem_20_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n13), .I3(GND_net), .O(n6239));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4766_3_lut (.I0(\REG.mem_20_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n13), .I3(GND_net), .O(n6240));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4767_3_lut (.I0(\REG.mem_20_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n13), .I3(GND_net), .O(n6241));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4768_3_lut (.I0(\REG.mem_20_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n13), .I3(GND_net), .O(n6242));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4769_3_lut (.I0(\REG.mem_20_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n13), .I3(GND_net), .O(n6243));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4770_3_lut (.I0(\REG.mem_20_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n13), .I3(GND_net), .O(n6244));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4770_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4771_3_lut (.I0(\REG.mem_20_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n13), .I3(GND_net), .O(n6245));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4772_3_lut (.I0(\REG.mem_20_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n13), .I3(GND_net), .O(n6246));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4773_3_lut (.I0(\REG.mem_20_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n13), .I3(GND_net), .O(n6247));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4774_3_lut (.I0(\REG.mem_20_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n13), .I3(GND_net), .O(n6248));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5476_3_lut (.I0(n5460), .I1(r_Bit_Index_adj_1469[0]), .I2(n5024), 
            .I3(GND_net), .O(n6950));   // src/uart_tx.v(38[10] 141[8])
    defparam i5476_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i4179_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[5]), .I2(\mem_LUT.data_raw_r [5]), 
            .I3(n5086), .O(n5653));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4179_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4174_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[6]), .I2(\mem_LUT.data_raw_r [6]), 
            .I3(n5086), .O(n5648));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4174_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4171_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[7]), .I2(\mem_LUT.data_raw_r [7]), 
            .I3(n5086), .O(n5645));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4171_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4775_3_lut (.I0(\REG.mem_20_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n13), .I3(GND_net), .O(n6249));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4776_3_lut (.I0(\REG.mem_20_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n13), .I3(GND_net), .O(n6250));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4777_3_lut (.I0(\REG.mem_20_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n13), .I3(GND_net), .O(n6251));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4778_3_lut (.I0(\REG.mem_20_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n13), .I3(GND_net), .O(n6252));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4779_3_lut (.I0(\REG.mem_20_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n13), .I3(GND_net), .O(n6253));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4780_3_lut (.I0(\REG.mem_20_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n13), .I3(GND_net), .O(n6254));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4781_3_lut (.I0(\REG.mem_20_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n13), .I3(GND_net), .O(n6255));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4782_3_lut (.I0(\REG.mem_20_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n13), .I3(GND_net), .O(n6256));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4783_3_lut (.I0(\REG.mem_20_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n13), .I3(GND_net), .O(n6257));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4784_3_lut (.I0(\REG.mem_20_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n13), .I3(GND_net), .O(n6258));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4785_3_lut (.I0(\REG.mem_20_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n13), .I3(GND_net), .O(n6259));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5482_3_lut (.I0(n13034), .I1(r_Bit_Index[0]), .I2(n13008), 
            .I3(GND_net), .O(n6956));   // src/uart_rx.v(49[10] 144[8])
    defparam i5482_3_lut.LUT_INIT = 16'h1414;
    \uart_rx(CLKS_PER_BIT=20)  pc_rx (.SLM_CLK_c(SLM_CLK_c), .r_Rx_Data(r_Rx_Data), 
            .r_Bit_Index({Open_0, Open_1, r_Bit_Index[0]}), .n4790(n4790), 
            .GND_net(GND_net), .n4(n4_adj_1435), .n6967(n6967), .pc_data_rx({pc_data_rx}), 
            .VCC_net(VCC_net), .debug_led3(debug_led3), .n6956(n6956), 
            .n6909(n6909), .n6908(n6908), .n6907(n6907), .n6906(n6906), 
            .n6905(n6905), .n6904(n6904), .n6903(n6903), .n13008(n13008), 
            .n13034(n13034), .UART_RX_c(UART_RX_c), .n4787(n4787), .n4_adj_9(n4_adj_1434), 
            .n4_adj_10(n4_adj_1436), .n4794(n4794)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(790[42] 795[3])
    SB_LUT4 i4786_3_lut (.I0(\REG.mem_20_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n13), .I3(GND_net), .O(n6260));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4973_3_lut (.I0(\REG.mem_26_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n7), .I3(GND_net), .O(n6447));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4161_2_lut (.I0(is_tx_fifo_full_flag), .I1(spi_rx_byte_ready), 
            .I2(GND_net), .I3(GND_net), .O(n5635));   // src/top.v(980[8] 989[4])
    defparam i4161_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4162_2_lut_3_lut (.I0(reset_all_w), .I1(fifo_read_cmd), .I2(is_fifo_empty_flag), 
            .I3(GND_net), .O(n5636));   // src/fifo_quad_word_mod.v(353[29] 363[32])
    defparam i4162_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i5467_3_lut_4_lut (.I0(r_SM_Main_2__N_1029[0]), .I1(fifo_read_cmd), 
            .I2(is_fifo_empty_flag), .I3(tx_uart_active_flag), .O(n6941));   // src/top.v(1001[8] 1019[4])
    defparam i5467_3_lut_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1114_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(n63), 
            .I3(state[2]), .O(n2335));   // src/timing_controller.v(78[11:16])
    defparam i1114_4_lut_4_lut.LUT_INIT = 16'h0806;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_1467[1]), .I1(r_SM_Main_2__N_1026[1]), 
            .I2(r_SM_Main_adj_1467[0]), .I3(r_SM_Main_adj_1467[2]), .O(n16231));   // src/uart_tx.v(38[10] 141[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0080;
    fifo_dc_32_lut_gen2 fifo_dc_32_lut_gen_inst (.dc32_fifo_data_in({dc32_fifo_data_in}), 
            .\REG.mem_1_9 (\REG.mem_1_9 ), .GND_net(GND_net), .\REG.mem_6_9 (\REG.mem_6_9 ), 
            .\REG.mem_7_9 (\REG.mem_7_9 ), .\REG.mem_4_9 (\REG.mem_4_9 ), 
            .\REG.mem_5_9 (\REG.mem_5_9 ), .\REG.mem_24_9 (\REG.mem_24_9 ), 
            .\REG.mem_25_9 (\REG.mem_25_9 ), .\REG.mem_1_31 (\REG.mem_1_31 ), 
            .\REG.mem_9_5 (\REG.mem_9_5 ), .\REG.mem_8_5 (\REG.mem_8_5 ), 
            .\REG.mem_26_9 (\REG.mem_26_9 ), .\REG.mem_27_9 (\REG.mem_27_9 ), 
            .rd_grey_sync_r({rd_grey_sync_r}), .\REG.mem_17_25 (\REG.mem_17_25 ), 
            .\REG.mem_6_16 (\REG.mem_6_16 ), .\REG.mem_7_16 (\REG.mem_7_16 ), 
            .\REG.mem_1_7 (\REG.mem_1_7 ), .\REG.mem_6_7 (\REG.mem_6_7 ), 
            .\REG.mem_7_7 (\REG.mem_7_7 ), .\REG.mem_4_7 (\REG.mem_4_7 ), 
            .\REG.mem_5_7 (\REG.mem_5_7 ), .\REG.mem_10_23 (\REG.mem_10_23 ), 
            .\REG.mem_11_23 (\REG.mem_11_23 ), .\REG.mem_5_16 (\REG.mem_5_16 ), 
            .\REG.mem_4_16 (\REG.mem_4_16 ), .\REG.mem_17_7 (\REG.mem_17_7 ), 
            .\REG.mem_22_7 (\REG.mem_22_7 ), .\REG.mem_23_7 (\REG.mem_23_7 ), 
            .\REG.mem_20_7 (\REG.mem_20_7 ), .\REG.mem_21_7 (\REG.mem_21_7 ), 
            .\REG.mem_9_23 (\REG.mem_9_23 ), .\REG.mem_8_23 (\REG.mem_8_23 ), 
            .n7(n7), .n23(n23), .FIFO_CLK_c(FIFO_CLK_c), .DEBUG_1_c(DEBUG_1_c), 
            .reset_per_frame(reset_per_frame), .wr_fifo_en_w(wr_fifo_en_w), 
            .\wr_addr_r[0] (wr_addr_r[0]), .\REG.mem_22_29 (\REG.mem_22_29 ), 
            .\REG.mem_23_29 (\REG.mem_23_29 ), .\REG.mem_21_29 (\REG.mem_21_29 ), 
            .\REG.mem_20_29 (\REG.mem_20_29 ), .DEBUG_5_c_0(DEBUG_5_c_0), 
            .SLM_CLK_c(SLM_CLK_c), .\REG.mem_26_21 (\REG.mem_26_21 ), .\REG.mem_27_21 (\REG.mem_27_21 ), 
            .\REG.mem_26_25 (\REG.mem_26_25 ), .\REG.mem_27_25 (\REG.mem_27_25 ), 
            .\REG.mem_25_25 (\REG.mem_25_25 ), .\REG.mem_24_25 (\REG.mem_24_25 ), 
            .\REG.mem_25_21 (\REG.mem_25_21 ), .\REG.mem_24_21 (\REG.mem_24_21 ), 
            .\REG.mem_1_10 (\REG.mem_1_10 ), .\REG.mem_6_10 (\REG.mem_6_10 ), 
            .\REG.mem_7_10 (\REG.mem_7_10 ), .\REG.mem_4_10 (\REG.mem_4_10 ), 
            .\REG.mem_5_10 (\REG.mem_5_10 ), .\REG.mem_1_26 (\REG.mem_1_26 ), 
            .n28(n28), .n12(n12), .dc32_fifo_empty(dc32_fifo_empty), .\wr_grey_sync_r[0] (wr_grey_sync_r[0]), 
            .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .dc32_fifo_almost_empty(dc32_fifo_almost_empty), .n32(n32), 
            .n16(n16), .\REG.mem_17_10 (\REG.mem_17_10 ), .\REG.mem_22_10 (\REG.mem_22_10 ), 
            .\REG.mem_23_10 (\REG.mem_23_10 ), .\REG.mem_20_10 (\REG.mem_20_10 ), 
            .\REG.mem_21_10 (\REG.mem_21_10 ), .dc32_fifo_full(dc32_fifo_full), 
            .\REG.mem_10_28 (\REG.mem_10_28 ), .\REG.mem_11_28 (\REG.mem_11_28 ), 
            .\REG.mem_9_28 (\REG.mem_9_28 ), .\REG.mem_8_28 (\REG.mem_8_28 ), 
            .\REG.mem_17_29 (\REG.mem_17_29 ), .\rd_addr_nxt_c_5__N_573[3] (rd_addr_nxt_c_5__N_573[3]), 
            .\rd_addr_nxt_c_5__N_573[1] (rd_addr_nxt_c_5__N_573[1]), .n6(n6), 
            .n22(n22), .\REG.mem_1_28 (\REG.mem_1_28 ), .\REG.mem_6_28 (\REG.mem_6_28 ), 
            .\REG.mem_7_28 (\REG.mem_7_28 ), .\REG.mem_4_28 (\REG.mem_4_28 ), 
            .\REG.mem_5_28 (\REG.mem_5_28 ), .\REG.mem_1_2 (\REG.mem_1_2 ), 
            .\REG.mem_6_2 (\REG.mem_6_2 ), .\REG.mem_7_2 (\REG.mem_7_2 ), 
            .\REG.mem_4_2 (\REG.mem_4_2 ), .\REG.mem_5_2 (\REG.mem_5_2 ), 
            .\REG.mem_1_22 (\REG.mem_1_22 ), .\REG.mem_6_22 (\REG.mem_6_22 ), 
            .\REG.mem_7_22 (\REG.mem_7_22 ), .\REG.mem_4_22 (\REG.mem_4_22 ), 
            .\REG.mem_5_22 (\REG.mem_5_22 ), .\REG.mem_17_22 (\REG.mem_17_22 ), 
            .\REG.mem_22_22 (\REG.mem_22_22 ), .\REG.mem_23_22 (\REG.mem_23_22 ), 
            .\REG.mem_20_22 (\REG.mem_20_22 ), .\REG.mem_21_22 (\REG.mem_21_22 ), 
            .\rd_addr_nxt_c_5__N_573[4] (rd_addr_nxt_c_5__N_573[4]), .\REG.mem_5_18 (\REG.mem_5_18 ), 
            .\REG.mem_4_18 (\REG.mem_4_18 ), .\REG.mem_6_4 (\REG.mem_6_4 ), 
            .\REG.mem_7_4 (\REG.mem_7_4 ), .\REG.mem_6_18 (\REG.mem_6_18 ), 
            .\REG.mem_7_18 (\REG.mem_7_18 ), .\REG.mem_10_8 (\REG.mem_10_8 ), 
            .\REG.mem_11_8 (\REG.mem_11_8 ), .\REG.mem_9_8 (\REG.mem_9_8 ), 
            .\REG.mem_8_8 (\REG.mem_8_8 ), .\REG.mem_5_4 (\REG.mem_5_4 ), 
            .\REG.mem_4_4 (\REG.mem_4_4 ), .\REG.mem_1_21 (\REG.mem_1_21 ), 
            .n7013(n7013), .n7012(n7012), .n7011(n7011), .n7010(n7010), 
            .n7009(n7009), .n7008(n7008), .wp_sync1_r({wp_sync1_r}), .n7007(n7007), 
            .n7006(n7006), .n7005(n7005), .n7004(n7004), .n7003(n7003), 
            .n7002(n7002), .n7000(n7000), .n6998(n6998), .n6997(n6997), 
            .n6996(n6996), .n6995(n6995), .n6994(n6994), .n6993(n6993), 
            .rp_sync1_r({rp_sync1_r}), .n6992(n6992), .n6991(n6991), .n6990(n6990), 
            .n6989(n6989), .\REG.mem_1_13 (\REG.mem_1_13 ), .n6930(n6930), 
            .n6928(n6928), .\wr_addr_r[5] (wr_addr_r[5]), .\REG.mem_6_30 (\REG.mem_6_30 ), 
            .\REG.mem_7_30 (\REG.mem_7_30 ), .n6493(n6493), .\REG.mem_27_31 (\REG.mem_27_31 ), 
            .n6492(n6492), .\REG.mem_27_30 (\REG.mem_27_30 ), .n6491(n6491), 
            .\REG.mem_27_29 (\REG.mem_27_29 ), .n6490(n6490), .\REG.mem_27_28 (\REG.mem_27_28 ), 
            .n6489(n6489), .\REG.mem_27_27 (\REG.mem_27_27 ), .n6488(n6488), 
            .\REG.mem_27_26 (\REG.mem_27_26 ), .n6487(n6487), .n6486(n6486), 
            .\REG.mem_27_24 (\REG.mem_27_24 ), .n6485(n6485), .\REG.mem_27_23 (\REG.mem_27_23 ), 
            .n6484(n6484), .\REG.mem_27_22 (\REG.mem_27_22 ), .n6483(n6483), 
            .n6482(n6482), .\REG.mem_27_20 (\REG.mem_27_20 ), .n6481(n6481), 
            .\REG.mem_27_19 (\REG.mem_27_19 ), .n6480(n6480), .\REG.mem_27_18 (\REG.mem_27_18 ), 
            .n6479(n6479), .\REG.mem_27_17 (\REG.mem_27_17 ), .n6478(n6478), 
            .\REG.mem_27_16 (\REG.mem_27_16 ), .n6477(n6477), .\REG.mem_27_15 (\REG.mem_27_15 ), 
            .n6476(n6476), .\REG.mem_27_14 (\REG.mem_27_14 ), .n6475(n6475), 
            .\REG.mem_27_13 (\REG.mem_27_13 ), .n6474(n6474), .\REG.mem_27_12 (\REG.mem_27_12 ), 
            .n6473(n6473), .\REG.mem_27_11 (\REG.mem_27_11 ), .n6472(n6472), 
            .\REG.mem_27_10 (\REG.mem_27_10 ), .n6471(n6471), .n6470(n6470), 
            .\REG.mem_27_8 (\REG.mem_27_8 ), .n6469(n6469), .\REG.mem_27_7 (\REG.mem_27_7 ), 
            .n6468(n6468), .\REG.mem_27_6 (\REG.mem_27_6 ), .n6467(n6467), 
            .\REG.mem_27_5 (\REG.mem_27_5 ), .n6466(n6466), .\REG.mem_27_4 (\REG.mem_27_4 ), 
            .n6465(n6465), .\REG.mem_27_3 (\REG.mem_27_3 ), .n6464(n6464), 
            .\REG.mem_27_2 (\REG.mem_27_2 ), .n6463(n6463), .\REG.mem_27_1 (\REG.mem_27_1 ), 
            .n6462(n6462), .\REG.mem_27_0 (\REG.mem_27_0 ), .n6461(n6461), 
            .\REG.mem_26_31 (\REG.mem_26_31 ), .n6460(n6460), .\REG.mem_26_30 (\REG.mem_26_30 ), 
            .n6459(n6459), .\REG.mem_26_29 (\REG.mem_26_29 ), .n6458(n6458), 
            .\REG.mem_26_28 (\REG.mem_26_28 ), .n6457(n6457), .\REG.mem_26_27 (\REG.mem_26_27 ), 
            .n6456(n6456), .\REG.mem_26_26 (\REG.mem_26_26 ), .n6455(n6455), 
            .n6454(n6454), .\REG.mem_26_24 (\REG.mem_26_24 ), .n6453(n6453), 
            .\REG.mem_26_23 (\REG.mem_26_23 ), .n6452(n6452), .\REG.mem_26_22 (\REG.mem_26_22 ), 
            .n6451(n6451), .n6450(n6450), .\REG.mem_26_20 (\REG.mem_26_20 ), 
            .n6449(n6449), .\REG.mem_26_19 (\REG.mem_26_19 ), .n6448(n6448), 
            .\REG.mem_26_18 (\REG.mem_26_18 ), .n6447(n6447), .\REG.mem_26_17 (\REG.mem_26_17 ), 
            .n6446(n6446), .\REG.mem_26_16 (\REG.mem_26_16 ), .n6445(n6445), 
            .\REG.mem_26_15 (\REG.mem_26_15 ), .n6444(n6444), .\REG.mem_26_14 (\REG.mem_26_14 ), 
            .n6443(n6443), .\REG.mem_26_13 (\REG.mem_26_13 ), .n6442(n6442), 
            .\REG.mem_26_12 (\REG.mem_26_12 ), .n6441(n6441), .\REG.mem_26_11 (\REG.mem_26_11 ), 
            .n6440(n6440), .\REG.mem_26_10 (\REG.mem_26_10 ), .n6439(n6439), 
            .n6438(n6438), .\REG.mem_26_8 (\REG.mem_26_8 ), .n6437(n6437), 
            .\REG.mem_26_7 (\REG.mem_26_7 ), .n6436(n6436), .\REG.mem_26_6 (\REG.mem_26_6 ), 
            .n6435(n6435), .\REG.mem_26_5 (\REG.mem_26_5 ), .n6434(n6434), 
            .\REG.mem_26_4 (\REG.mem_26_4 ), .n6433(n6433), .\REG.mem_26_3 (\REG.mem_26_3 ), 
            .n6432(n6432), .\REG.mem_26_2 (\REG.mem_26_2 ), .n6431(n6431), 
            .\REG.mem_26_1 (\REG.mem_26_1 ), .n6430(n6430), .\REG.mem_26_0 (\REG.mem_26_0 ), 
            .n6429(n6429), .\REG.mem_25_31 (\REG.mem_25_31 ), .n6428(n6428), 
            .\REG.mem_25_30 (\REG.mem_25_30 ), .n6427(n6427), .\REG.mem_25_29 (\REG.mem_25_29 ), 
            .n6426(n6426), .\REG.mem_25_28 (\REG.mem_25_28 ), .n6425(n6425), 
            .\REG.mem_25_27 (\REG.mem_25_27 ), .n6424(n6424), .\REG.mem_25_26 (\REG.mem_25_26 ), 
            .n6423(n6423), .n6422(n6422), .\REG.mem_25_24 (\REG.mem_25_24 ), 
            .n6421(n6421), .\REG.mem_25_23 (\REG.mem_25_23 ), .n6420(n6420), 
            .\REG.mem_25_22 (\REG.mem_25_22 ), .n6419(n6419), .n6418(n6418), 
            .\REG.mem_25_20 (\REG.mem_25_20 ), .n6417(n6417), .\REG.mem_25_19 (\REG.mem_25_19 ), 
            .n6416(n6416), .\REG.mem_25_18 (\REG.mem_25_18 ), .n6415(n6415), 
            .\REG.mem_25_17 (\REG.mem_25_17 ), .n6414(n6414), .\REG.mem_25_16 (\REG.mem_25_16 ), 
            .n6413(n6413), .\REG.mem_25_15 (\REG.mem_25_15 ), .n6412(n6412), 
            .\REG.mem_25_14 (\REG.mem_25_14 ), .n6411(n6411), .\REG.mem_25_13 (\REG.mem_25_13 ), 
            .n6410(n6410), .\REG.mem_25_12 (\REG.mem_25_12 ), .n6409(n6409), 
            .\REG.mem_25_11 (\REG.mem_25_11 ), .n6408(n6408), .\REG.mem_25_10 (\REG.mem_25_10 ), 
            .n6407(n6407), .n6406(n6406), .\REG.mem_25_8 (\REG.mem_25_8 ), 
            .n6405(n6405), .\REG.mem_25_7 (\REG.mem_25_7 ), .n6404(n6404), 
            .\REG.mem_25_6 (\REG.mem_25_6 ), .n6403(n6403), .\REG.mem_25_5 (\REG.mem_25_5 ), 
            .n6402(n6402), .\REG.mem_25_4 (\REG.mem_25_4 ), .n6401(n6401), 
            .\REG.mem_25_3 (\REG.mem_25_3 ), .n6400(n6400), .\REG.mem_25_2 (\REG.mem_25_2 ), 
            .n6399(n6399), .\REG.mem_25_1 (\REG.mem_25_1 ), .n6398(n6398), 
            .\REG.mem_25_0 (\REG.mem_25_0 ), .n6397(n6397), .\REG.mem_24_31 (\REG.mem_24_31 ), 
            .n6396(n6396), .\REG.mem_24_30 (\REG.mem_24_30 ), .n6395(n6395), 
            .\REG.mem_24_29 (\REG.mem_24_29 ), .n6394(n6394), .\REG.mem_24_28 (\REG.mem_24_28 ), 
            .n6393(n6393), .\REG.mem_24_27 (\REG.mem_24_27 ), .n6392(n6392), 
            .\REG.mem_24_26 (\REG.mem_24_26 ), .n6391(n6391), .n6390(n6390), 
            .\REG.mem_24_24 (\REG.mem_24_24 ), .n6389(n6389), .\REG.mem_24_23 (\REG.mem_24_23 ), 
            .n6388(n6388), .\REG.mem_24_22 (\REG.mem_24_22 ), .n6387(n6387), 
            .n6386(n6386), .\REG.mem_24_20 (\REG.mem_24_20 ), .n6385(n6385), 
            .\REG.mem_24_19 (\REG.mem_24_19 ), .n6384(n6384), .\REG.mem_24_18 (\REG.mem_24_18 ), 
            .n6383(n6383), .\REG.mem_24_17 (\REG.mem_24_17 ), .n6382(n6382), 
            .\REG.mem_24_16 (\REG.mem_24_16 ), .n6381(n6381), .\REG.mem_24_15 (\REG.mem_24_15 ), 
            .n6380(n6380), .\REG.mem_24_14 (\REG.mem_24_14 ), .n6379(n6379), 
            .\REG.mem_24_13 (\REG.mem_24_13 ), .n6378(n6378), .\REG.mem_24_12 (\REG.mem_24_12 ), 
            .n6377(n6377), .\REG.mem_24_11 (\REG.mem_24_11 ), .n6376(n6376), 
            .\REG.mem_24_10 (\REG.mem_24_10 ), .n6375(n6375), .n6374(n6374), 
            .\REG.mem_24_8 (\REG.mem_24_8 ), .n6373(n6373), .\REG.mem_24_7 (\REG.mem_24_7 ), 
            .n6372(n6372), .\REG.mem_24_6 (\REG.mem_24_6 ), .n6371(n6371), 
            .\REG.mem_24_5 (\REG.mem_24_5 ), .n6370(n6370), .\REG.mem_24_4 (\REG.mem_24_4 ), 
            .n6369(n6369), .\REG.mem_24_3 (\REG.mem_24_3 ), .n6368(n6368), 
            .\REG.mem_24_2 (\REG.mem_24_2 ), .n6367(n6367), .\REG.mem_24_1 (\REG.mem_24_1 ), 
            .n6366(n6366), .\REG.mem_24_0 (\REG.mem_24_0 ), .n6365(n6365), 
            .\REG.mem_23_31 (\REG.mem_23_31 ), .n6364(n6364), .\REG.mem_23_30 (\REG.mem_23_30 ), 
            .n6363(n6363), .n6362(n6362), .\REG.mem_23_28 (\REG.mem_23_28 ), 
            .n6361(n6361), .\REG.mem_23_27 (\REG.mem_23_27 ), .n6360(n6360), 
            .\REG.mem_23_26 (\REG.mem_23_26 ), .n6359(n6359), .\REG.mem_23_25 (\REG.mem_23_25 ), 
            .n6358(n6358), .\REG.mem_23_24 (\REG.mem_23_24 ), .n6357(n6357), 
            .\REG.mem_23_23 (\REG.mem_23_23 ), .n6356(n6356), .n6355(n6355), 
            .\REG.mem_23_21 (\REG.mem_23_21 ), .n6354(n6354), .\REG.mem_23_20 (\REG.mem_23_20 ), 
            .n6353(n6353), .\REG.mem_23_19 (\REG.mem_23_19 ), .n6352(n6352), 
            .\REG.mem_23_18 (\REG.mem_23_18 ), .n6351(n6351), .\REG.mem_23_17 (\REG.mem_23_17 ), 
            .n6350(n6350), .\REG.mem_23_16 (\REG.mem_23_16 ), .n6349(n6349), 
            .\REG.mem_23_15 (\REG.mem_23_15 ), .n6348(n6348), .\REG.mem_23_14 (\REG.mem_23_14 ), 
            .n6347(n6347), .\REG.mem_23_13 (\REG.mem_23_13 ), .n6346(n6346), 
            .\REG.mem_23_12 (\REG.mem_23_12 ), .n6345(n6345), .\REG.mem_23_11 (\REG.mem_23_11 ), 
            .n6344(n6344), .n6343(n6343), .\REG.mem_23_9 (\REG.mem_23_9 ), 
            .n6342(n6342), .\REG.mem_23_8 (\REG.mem_23_8 ), .n6341(n6341), 
            .n6340(n6340), .\REG.mem_23_6 (\REG.mem_23_6 ), .n6339(n6339), 
            .\REG.mem_23_5 (\REG.mem_23_5 ), .n6338(n6338), .\REG.mem_23_4 (\REG.mem_23_4 ), 
            .n6337(n6337), .\REG.mem_23_3 (\REG.mem_23_3 ), .n6336(n6336), 
            .\REG.mem_23_2 (\REG.mem_23_2 ), .n6335(n6335), .\REG.mem_23_1 (\REG.mem_23_1 ), 
            .n6334(n6334), .\REG.mem_23_0 (\REG.mem_23_0 ), .n6333(n6333), 
            .\REG.mem_22_31 (\REG.mem_22_31 ), .n6332(n6332), .\REG.mem_22_30 (\REG.mem_22_30 ), 
            .n6331(n6331), .n6330(n6330), .\REG.mem_22_28 (\REG.mem_22_28 ), 
            .n6329(n6329), .\REG.mem_22_27 (\REG.mem_22_27 ), .n6328(n6328), 
            .\REG.mem_22_26 (\REG.mem_22_26 ), .n6327(n6327), .\REG.mem_22_25 (\REG.mem_22_25 ), 
            .n6326(n6326), .\REG.mem_22_24 (\REG.mem_22_24 ), .n6325(n6325), 
            .\REG.mem_22_23 (\REG.mem_22_23 ), .n6324(n6324), .n6323(n6323), 
            .\REG.mem_22_21 (\REG.mem_22_21 ), .n6322(n6322), .\REG.mem_22_20 (\REG.mem_22_20 ), 
            .n6321(n6321), .\REG.mem_22_19 (\REG.mem_22_19 ), .n6320(n6320), 
            .\REG.mem_22_18 (\REG.mem_22_18 ), .n6319(n6319), .\REG.mem_22_17 (\REG.mem_22_17 ), 
            .n6318(n6318), .\REG.mem_22_16 (\REG.mem_22_16 ), .n6317(n6317), 
            .\REG.mem_22_15 (\REG.mem_22_15 ), .n6316(n6316), .\REG.mem_22_14 (\REG.mem_22_14 ), 
            .n6315(n6315), .\REG.mem_22_13 (\REG.mem_22_13 ), .n6314(n6314), 
            .\REG.mem_22_12 (\REG.mem_22_12 ), .n6313(n6313), .\REG.mem_22_11 (\REG.mem_22_11 ), 
            .n6312(n6312), .n6311(n6311), .\REG.mem_22_9 (\REG.mem_22_9 ), 
            .n6310(n6310), .\REG.mem_22_8 (\REG.mem_22_8 ), .n6309(n6309), 
            .n6308(n6308), .\REG.mem_22_6 (\REG.mem_22_6 ), .n6307(n6307), 
            .\REG.mem_22_5 (\REG.mem_22_5 ), .n6306(n6306), .\REG.mem_22_4 (\REG.mem_22_4 ), 
            .n6305(n6305), .\REG.mem_22_3 (\REG.mem_22_3 ), .n6304(n6304), 
            .\REG.mem_22_2 (\REG.mem_22_2 ), .n6303(n6303), .\REG.mem_22_1 (\REG.mem_22_1 ), 
            .n6302(n6302), .\REG.mem_22_0 (\REG.mem_22_0 ), .n6301(n6301), 
            .\REG.mem_21_31 (\REG.mem_21_31 ), .n6300(n6300), .\REG.mem_21_30 (\REG.mem_21_30 ), 
            .n6299(n6299), .n6298(n6298), .\REG.mem_21_28 (\REG.mem_21_28 ), 
            .n6297(n6297), .\REG.mem_21_27 (\REG.mem_21_27 ), .n6296(n6296), 
            .\REG.mem_21_26 (\REG.mem_21_26 ), .n6295(n6295), .\REG.mem_21_25 (\REG.mem_21_25 ), 
            .n6294(n6294), .\REG.mem_21_24 (\REG.mem_21_24 ), .n6293(n6293), 
            .\REG.mem_21_23 (\REG.mem_21_23 ), .n6292(n6292), .n6291(n6291), 
            .\REG.mem_21_21 (\REG.mem_21_21 ), .n6290(n6290), .\REG.mem_21_20 (\REG.mem_21_20 ), 
            .n6289(n6289), .\REG.mem_21_19 (\REG.mem_21_19 ), .n6288(n6288), 
            .\REG.mem_21_18 (\REG.mem_21_18 ), .n6287(n6287), .\REG.mem_21_17 (\REG.mem_21_17 ), 
            .n6286(n6286), .\REG.mem_21_16 (\REG.mem_21_16 ), .n6285(n6285), 
            .\REG.mem_21_15 (\REG.mem_21_15 ), .n6284(n6284), .\REG.mem_21_14 (\REG.mem_21_14 ), 
            .n6283(n6283), .\REG.mem_21_13 (\REG.mem_21_13 ), .n6282(n6282), 
            .\REG.mem_21_12 (\REG.mem_21_12 ), .n6281(n6281), .\REG.mem_21_11 (\REG.mem_21_11 ), 
            .n6280(n6280), .n6279(n6279), .\REG.mem_21_9 (\REG.mem_21_9 ), 
            .n6278(n6278), .\REG.mem_21_8 (\REG.mem_21_8 ), .n6277(n6277), 
            .n6276(n6276), .\REG.mem_21_6 (\REG.mem_21_6 ), .n6275(n6275), 
            .\REG.mem_21_5 (\REG.mem_21_5 ), .n6274(n6274), .\REG.mem_21_4 (\REG.mem_21_4 ), 
            .n6273(n6273), .\REG.mem_21_3 (\REG.mem_21_3 ), .n6272(n6272), 
            .\REG.mem_21_2 (\REG.mem_21_2 ), .n6271(n6271), .\REG.mem_21_1 (\REG.mem_21_1 ), 
            .n6270(n6270), .\REG.mem_21_0 (\REG.mem_21_0 ), .n6269(n6269), 
            .\REG.mem_20_31 (\REG.mem_20_31 ), .n6268(n6268), .\REG.mem_20_30 (\REG.mem_20_30 ), 
            .n6267(n6267), .n6266(n6266), .\REG.mem_20_28 (\REG.mem_20_28 ), 
            .n6265(n6265), .\REG.mem_20_27 (\REG.mem_20_27 ), .n6264(n6264), 
            .\REG.mem_20_26 (\REG.mem_20_26 ), .n6263(n6263), .\REG.mem_20_25 (\REG.mem_20_25 ), 
            .n6262(n6262), .\REG.mem_20_24 (\REG.mem_20_24 ), .n6261(n6261), 
            .\REG.mem_20_23 (\REG.mem_20_23 ), .n6260(n6260), .n6259(n6259), 
            .\REG.mem_20_21 (\REG.mem_20_21 ), .n6258(n6258), .\REG.mem_20_20 (\REG.mem_20_20 ), 
            .n6257(n6257), .\REG.mem_20_19 (\REG.mem_20_19 ), .n6256(n6256), 
            .\REG.mem_20_18 (\REG.mem_20_18 ), .n6255(n6255), .\REG.mem_20_17 (\REG.mem_20_17 ), 
            .n6254(n6254), .\REG.mem_20_16 (\REG.mem_20_16 ), .n6253(n6253), 
            .\REG.mem_20_15 (\REG.mem_20_15 ), .n6252(n6252), .\REG.mem_20_14 (\REG.mem_20_14 ), 
            .n6251(n6251), .\REG.mem_20_13 (\REG.mem_20_13 ), .n6250(n6250), 
            .\REG.mem_20_12 (\REG.mem_20_12 ), .n6249(n6249), .\REG.mem_20_11 (\REG.mem_20_11 ), 
            .n6248(n6248), .n6247(n6247), .\REG.mem_20_9 (\REG.mem_20_9 ), 
            .n6246(n6246), .\REG.mem_20_8 (\REG.mem_20_8 ), .n6245(n6245), 
            .n6244(n6244), .\REG.mem_20_6 (\REG.mem_20_6 ), .n6243(n6243), 
            .\REG.mem_20_5 (\REG.mem_20_5 ), .n6242(n6242), .\REG.mem_20_4 (\REG.mem_20_4 ), 
            .n6241(n6241), .\REG.mem_20_3 (\REG.mem_20_3 ), .n6240(n6240), 
            .\REG.mem_20_2 (\REG.mem_20_2 ), .n6239(n6239), .\REG.mem_20_1 (\REG.mem_20_1 ), 
            .n6238(n6238), .\REG.mem_20_0 (\REG.mem_20_0 ), .n6173(n6173), 
            .\REG.mem_17_31 (\REG.mem_17_31 ), .n6172(n6172), .\REG.mem_17_30 (\REG.mem_17_30 ), 
            .n6171(n6171), .n6170(n6170), .\REG.mem_17_28 (\REG.mem_17_28 ), 
            .n6169(n6169), .\REG.mem_17_27 (\REG.mem_17_27 ), .n6168(n6168), 
            .\REG.mem_17_26 (\REG.mem_17_26 ), .n6167(n6167), .n6166(n6166), 
            .\REG.mem_17_24 (\REG.mem_17_24 ), .n6165(n6165), .\REG.mem_17_23 (\REG.mem_17_23 ), 
            .n6164(n6164), .n6163(n6163), .\REG.mem_17_21 (\REG.mem_17_21 ), 
            .n6162(n6162), .\REG.mem_17_20 (\REG.mem_17_20 ), .n6161(n6161), 
            .\REG.mem_17_19 (\REG.mem_17_19 ), .n6160(n6160), .\REG.mem_17_18 (\REG.mem_17_18 ), 
            .n6159(n6159), .\REG.mem_17_17 (\REG.mem_17_17 ), .n6158(n6158), 
            .\REG.mem_17_16 (\REG.mem_17_16 ), .n6157(n6157), .\REG.mem_17_15 (\REG.mem_17_15 ), 
            .n6156(n6156), .\REG.mem_17_14 (\REG.mem_17_14 ), .n6155(n6155), 
            .\REG.mem_17_13 (\REG.mem_17_13 ), .n6154(n6154), .\REG.mem_17_12 (\REG.mem_17_12 ), 
            .n6153(n6153), .\REG.mem_17_11 (\REG.mem_17_11 ), .n6152(n6152), 
            .n6151(n6151), .\REG.mem_17_9 (\REG.mem_17_9 ), .n6150(n6150), 
            .\REG.mem_17_8 (\REG.mem_17_8 ), .n6149(n6149), .n6148(n6148), 
            .\REG.mem_17_6 (\REG.mem_17_6 ), .n6147(n6147), .\REG.mem_17_5 (\REG.mem_17_5 ), 
            .n6146(n6146), .\REG.mem_17_4 (\REG.mem_17_4 ), .n6145(n6145), 
            .\REG.mem_17_3 (\REG.mem_17_3 ), .n6144(n6144), .\REG.mem_17_2 (\REG.mem_17_2 ), 
            .n6143(n6143), .\REG.mem_17_1 (\REG.mem_17_1 ), .n6142(n6142), 
            .\REG.mem_17_0 (\REG.mem_17_0 ), .\REG.mem_5_30 (\REG.mem_5_30 ), 
            .\REG.mem_4_30 (\REG.mem_4_30 ), .\REG.mem_1_1 (\REG.mem_1_1 ), 
            .\REG.mem_6_1 (\REG.mem_6_1 ), .\REG.mem_7_1 (\REG.mem_7_1 ), 
            .\REG.mem_4_1 (\REG.mem_4_1 ), .\REG.mem_5_1 (\REG.mem_5_1 ), 
            .\REG.mem_6_21 (\REG.mem_6_21 ), .\REG.mem_7_21 (\REG.mem_7_21 ), 
            .\REG.mem_5_21 (\REG.mem_5_21 ), .\REG.mem_4_21 (\REG.mem_4_21 ), 
            .\REG.mem_1_30 (\REG.mem_1_30 ), .\REG.mem_10_21 (\REG.mem_10_21 ), 
            .\REG.mem_11_21 (\REG.mem_11_21 ), .\REG.mem_1_19 (\REG.mem_1_19 ), 
            .\REG.mem_6_19 (\REG.mem_6_19 ), .\REG.mem_7_19 (\REG.mem_7_19 ), 
            .\REG.mem_5_19 (\REG.mem_5_19 ), .\REG.mem_4_19 (\REG.mem_4_19 ), 
            .\REG.mem_9_21 (\REG.mem_9_21 ), .\REG.mem_8_21 (\REG.mem_8_21 ), 
            .\wr_addr_p1_w[0] (wr_addr_p1_w[0]), .\REG.mem_6_13 (\REG.mem_6_13 ), 
            .\REG.mem_7_13 (\REG.mem_7_13 ), .\REG.mem_5_13 (\REG.mem_5_13 ), 
            .\REG.mem_4_13 (\REG.mem_4_13 ), .\REG.mem_10_13 (\REG.mem_10_13 ), 
            .\REG.mem_11_13 (\REG.mem_11_13 ), .\REG.mem_9_13 (\REG.mem_9_13 ), 
            .\REG.mem_8_13 (\REG.mem_8_13 ), .\REG.mem_10_19 (\REG.mem_10_19 ), 
            .\REG.mem_11_19 (\REG.mem_11_19 ), .\REG.mem_9_19 (\REG.mem_9_19 ), 
            .\REG.mem_8_19 (\REG.mem_8_19 ), .\REG.mem_1_27 (\REG.mem_1_27 ), 
            .\REG.mem_6_27 (\REG.mem_6_27 ), .\REG.mem_7_27 (\REG.mem_7_27 ), 
            .\REG.mem_4_27 (\REG.mem_4_27 ), .\REG.mem_5_27 (\REG.mem_5_27 ), 
            .\REG.mem_1_6 (\REG.mem_1_6 ), .\REG.mem_8_2 (\REG.mem_8_2 ), 
            .\REG.mem_9_2 (\REG.mem_9_2 ), .\REG.mem_10_2 (\REG.mem_10_2 ), 
            .\REG.mem_11_2 (\REG.mem_11_2 ), .\wr_addr_nxt_c[2] (wr_addr_nxt_c[2]), 
            .VCC_net(VCC_net), .dc32_fifo_write_enable(dc32_fifo_write_enable), 
            .\REG.mem_1_0 (\REG.mem_1_0 ), .\REG.mem_10_15 (\REG.mem_10_15 ), 
            .\REG.mem_11_15 (\REG.mem_11_15 ), .\REG.mem_9_15 (\REG.mem_9_15 ), 
            .\REG.mem_8_15 (\REG.mem_8_15 ), .\dc32_fifo_data_out[1] (dc32_fifo_data_out[1]), 
            .\REG.mem_10_11 (\REG.mem_10_11 ), .\REG.mem_11_11 (\REG.mem_11_11 ), 
            .\REG.mem_9_11 (\REG.mem_9_11 ), .\REG.mem_8_11 (\REG.mem_8_11 ), 
            .\dc32_fifo_data_out[2] (dc32_fifo_data_out[2]), .\dc32_fifo_data_out[3] (dc32_fifo_data_out[3]), 
            .\dc32_fifo_data_out[4] (dc32_fifo_data_out[4]), .\dc32_fifo_data_out[5] (dc32_fifo_data_out[5]), 
            .\dc32_fifo_data_out[6] (dc32_fifo_data_out[6]), .\dc32_fifo_data_out[7] (dc32_fifo_data_out[7]), 
            .\dc32_fifo_data_out[8] (dc32_fifo_data_out[8]), .\dc32_fifo_data_out[9] (dc32_fifo_data_out[9]), 
            .\dc32_fifo_data_out[10] (dc32_fifo_data_out[10]), .\dc32_fifo_data_out[11] (dc32_fifo_data_out[11]), 
            .\dc32_fifo_data_out[12] (dc32_fifo_data_out[12]), .\dc32_fifo_data_out[13] (dc32_fifo_data_out[13]), 
            .\dc32_fifo_data_out[14] (dc32_fifo_data_out[14]), .\dc32_fifo_data_out[15] (dc32_fifo_data_out[15]), 
            .\dc32_fifo_data_out[16] (dc32_fifo_data_out[16]), .\dc32_fifo_data_out[17] (dc32_fifo_data_out[17]), 
            .\dc32_fifo_data_out[18] (dc32_fifo_data_out[18]), .\dc32_fifo_data_out[19] (dc32_fifo_data_out[19]), 
            .\dc32_fifo_data_out[20] (dc32_fifo_data_out[20]), .\dc32_fifo_data_out[21] (dc32_fifo_data_out[21]), 
            .\dc32_fifo_data_out[22] (dc32_fifo_data_out[22]), .\dc32_fifo_data_out[23] (dc32_fifo_data_out[23]), 
            .\dc32_fifo_data_out[24] (dc32_fifo_data_out[24]), .\dc32_fifo_data_out[25] (dc32_fifo_data_out[25]), 
            .\dc32_fifo_data_out[26] (dc32_fifo_data_out[26]), .\dc32_fifo_data_out[27] (dc32_fifo_data_out[27]), 
            .\dc32_fifo_data_out[28] (dc32_fifo_data_out[28]), .\dc32_fifo_data_out[29] (dc32_fifo_data_out[29]), 
            .\dc32_fifo_data_out[30] (dc32_fifo_data_out[30]), .\dc32_fifo_data_out[31] (dc32_fifo_data_out[31]), 
            .n7_adj_6(n7_adj_1420), .n8(n8_adj_1439), .n25(n25_adj_1444), 
            .n5981(n5981), .\REG.mem_11_31 (\REG.mem_11_31 ), .\REG.mem_1_23 (\REG.mem_1_23 ), 
            .n5980(n5980), .\REG.mem_11_30 (\REG.mem_11_30 ), .\REG.mem_6_6 (\REG.mem_6_6 ), 
            .\REG.mem_7_6 (\REG.mem_7_6 ), .\REG.mem_5_6 (\REG.mem_5_6 ), 
            .\REG.mem_4_6 (\REG.mem_4_6 ), .n5979(n5979), .\REG.mem_11_29 (\REG.mem_11_29 ), 
            .\REG.mem_10_29 (\REG.mem_10_29 ), .n5978(n5978), .n5977(n5977), 
            .\REG.mem_11_27 (\REG.mem_11_27 ), .n5976(n5976), .\REG.mem_11_26 (\REG.mem_11_26 ), 
            .n5975(n5975), .\REG.mem_11_25 (\REG.mem_11_25 ), .n5974(n5974), 
            .\REG.mem_11_24 (\REG.mem_11_24 ), .\REG.mem_9_29 (\REG.mem_9_29 ), 
            .\REG.mem_8_29 (\REG.mem_8_29 ), .n5973(n5973), .n5972(n5972), 
            .\REG.mem_11_22 (\REG.mem_11_22 ), .n29(n29), .\REG.mem_8_17 (\REG.mem_8_17 ), 
            .\REG.mem_9_17 (\REG.mem_9_17 ), .\REG.mem_10_17 (\REG.mem_10_17 ), 
            .\REG.mem_11_17 (\REG.mem_11_17 ), .\REG.mem_1_24 (\REG.mem_1_24 ), 
            .n5971(n5971), .n5970(n5970), .\REG.mem_11_20 (\REG.mem_11_20 ), 
            .\REG.mem_6_31 (\REG.mem_6_31 ), .\REG.mem_7_31 (\REG.mem_7_31 ), 
            .\REG.mem_5_31 (\REG.mem_5_31 ), .\REG.mem_4_31 (\REG.mem_4_31 ), 
            .\wr_grey_sync_r[1] (wr_grey_sync_r[1]), .n24(n24), .n13(n13), 
            .n8_adj_7(n8_adj_1419), .\REG.mem_6_23 (\REG.mem_6_23 ), .\REG.mem_7_23 (\REG.mem_7_23 ), 
            .\REG.mem_5_23 (\REG.mem_5_23 ), .\REG.mem_4_23 (\REG.mem_4_23 ), 
            .\REG.mem_10_6 (\REG.mem_10_6 ), .\REG.mem_11_6 (\REG.mem_11_6 ), 
            .n5969(n5969), .\REG.mem_9_6 (\REG.mem_9_6 ), .\REG.mem_8_6 (\REG.mem_8_6 ), 
            .\wr_grey_sync_r[2] (wr_grey_sync_r[2]), .\wr_grey_sync_r[3] (wr_grey_sync_r[3]), 
            .\wr_grey_sync_r[4] (wr_grey_sync_r[4]), .n5968(n5968), .\REG.mem_11_18 (\REG.mem_11_18 ), 
            .n5967(n5967), .n5966(n5966), .\REG.mem_11_16 (\REG.mem_11_16 ), 
            .n5965(n5965), .n5964(n5964), .\REG.mem_11_14 (\REG.mem_11_14 ), 
            .n5963(n5963), .n5962(n5962), .\REG.mem_11_12 (\REG.mem_11_12 ), 
            .n5961(n5961), .n5960(n5960), .\REG.mem_11_10 (\REG.mem_11_10 ), 
            .n5959(n5959), .\REG.mem_11_9 (\REG.mem_11_9 ), .n5958(n5958), 
            .n5957(n5957), .\REG.mem_11_7 (\REG.mem_11_7 ), .n5956(n5956), 
            .n5955(n5955), .\REG.mem_11_5 (\REG.mem_11_5 ), .n5954(n5954), 
            .\REG.mem_11_4 (\REG.mem_11_4 ), .n5953(n5953), .\REG.mem_11_3 (\REG.mem_11_3 ), 
            .\REG.mem_10_22 (\REG.mem_10_22 ), .n5952(n5952), .n5951(n5951), 
            .\REG.mem_11_1 (\REG.mem_11_1 ), .n5950(n5950), .\REG.mem_11_0 (\REG.mem_11_0 ), 
            .n5949(n5949), .\REG.mem_10_31 (\REG.mem_10_31 ), .n5948(n5948), 
            .\REG.mem_10_30 (\REG.mem_10_30 ), .n5947(n5947), .n5946(n5946), 
            .n5945(n5945), .\REG.mem_10_27 (\REG.mem_10_27 ), .\REG.mem_9_22 (\REG.mem_9_22 ), 
            .\REG.mem_8_22 (\REG.mem_8_22 ), .n5944(n5944), .\REG.mem_10_26 (\REG.mem_10_26 ), 
            .\REG.mem_1_18 (\REG.mem_1_18 ), .n5943(n5943), .\REG.mem_10_25 (\REG.mem_10_25 ), 
            .n5942(n5942), .\REG.mem_10_24 (\REG.mem_10_24 ), .n5611(n5611), 
            .\REG.mem_6_24 (\REG.mem_6_24 ), .\REG.mem_7_24 (\REG.mem_7_24 ), 
            .\REG.mem_5_24 (\REG.mem_5_24 ), .\REG.mem_4_24 (\REG.mem_4_24 ), 
            .\REG.mem_1_4 (\REG.mem_1_4 ), .\REG.mem_9_24 (\REG.mem_9_24 ), 
            .\REG.mem_8_24 (\REG.mem_8_24 ), .\REG.mem_6_0 (\REG.mem_6_0 ), 
            .\REG.mem_7_0 (\REG.mem_7_0 ), .\REG.mem_5_0 (\REG.mem_5_0 ), 
            .\REG.mem_4_0 (\REG.mem_4_0 ), .\REG.mem_10_4 (\REG.mem_10_4 ), 
            .n5610(n5610), .n5941(n5941), .n5940(n5940), .n5939(n5939), 
            .n5938(n5938), .\REG.mem_10_20 (\REG.mem_10_20 ), .n5937(n5937), 
            .n5608(n5608), .n5604(n5604), .n5603(n5603), .n5602(n5602), 
            .n5936(n5936), .\REG.mem_10_18 (\REG.mem_10_18 ), .n5935(n5935), 
            .n5934(n5934), .\REG.mem_10_16 (\REG.mem_10_16 ), .n5933(n5933), 
            .\REG.mem_1_17 (\REG.mem_1_17 ), .\REG.mem_9_4 (\REG.mem_9_4 ), 
            .\REG.mem_8_4 (\REG.mem_8_4 ), .\REG.mem_6_17 (\REG.mem_6_17 ), 
            .\REG.mem_7_17 (\REG.mem_7_17 ), .\REG.mem_4_17 (\REG.mem_4_17 ), 
            .\REG.mem_5_17 (\REG.mem_5_17 ), .dc32_fifo_read_enable(dc32_fifo_read_enable), 
            .n5932(n5932), .\REG.mem_10_14 (\REG.mem_10_14 ), .n5931(n5931), 
            .n5930(n5930), .\REG.mem_10_12 (\REG.mem_10_12 ), .n5929(n5929), 
            .n5928(n5928), .\REG.mem_10_10 (\REG.mem_10_10 ), .n5927(n5927), 
            .\REG.mem_10_9 (\REG.mem_10_9 ), .n5926(n5926), .n5925(n5925), 
            .\REG.mem_10_7 (\REG.mem_10_7 ), .n5924(n5924), .n5923(n5923), 
            .\REG.mem_10_5 (\REG.mem_10_5 ), .n5922(n5922), .n5921(n5921), 
            .\REG.mem_10_3 (\REG.mem_10_3 ), .n5920(n5920), .n5919(n5919), 
            .\REG.mem_10_1 (\REG.mem_10_1 ), .n5918(n5918), .\REG.mem_10_0 (\REG.mem_10_0 ), 
            .n5917(n5917), .\REG.mem_9_31 (\REG.mem_9_31 ), .n5916(n5916), 
            .\REG.mem_9_30 (\REG.mem_9_30 ), .n5915(n5915), .n5914(n5914), 
            .n5913(n5913), .\REG.mem_9_27 (\REG.mem_9_27 ), .n5912(n5912), 
            .\REG.mem_9_26 (\REG.mem_9_26 ), .n5911(n5911), .\REG.mem_9_25 (\REG.mem_9_25 ), 
            .n5910(n5910), .n5909(n5909), .n5908(n5908), .n5907(n5907), 
            .n5906(n5906), .\REG.mem_9_20 (\REG.mem_9_20 ), .n5905(n5905), 
            .n5904(n5904), .\REG.mem_9_18 (\REG.mem_9_18 ), .n5903(n5903), 
            .n5902(n5902), .\REG.mem_9_16 (\REG.mem_9_16 ), .n5901(n5901), 
            .n5900(n5900), .\REG.mem_9_14 (\REG.mem_9_14 ), .n5899(n5899), 
            .n5898(n5898), .\REG.mem_9_12 (\REG.mem_9_12 ), .n5897(n5897), 
            .n5896(n5896), .\REG.mem_9_10 (\REG.mem_9_10 ), .n5895(n5895), 
            .\REG.mem_9_9 (\REG.mem_9_9 ), .n5894(n5894), .n5893(n5893), 
            .\REG.mem_9_7 (\REG.mem_9_7 ), .n5892(n5892), .n5891(n5891), 
            .n5890(n5890), .n5889(n5889), .\REG.mem_9_3 (\REG.mem_9_3 ), 
            .n5888(n5888), .n5887(n5887), .\REG.mem_9_1 (\REG.mem_9_1 ), 
            .n5886(n5886), .\REG.mem_9_0 (\REG.mem_9_0 ), .n5885(n5885), 
            .\REG.mem_8_31 (\REG.mem_8_31 ), .n5884(n5884), .\REG.mem_8_30 (\REG.mem_8_30 ), 
            .n5883(n5883), .n5882(n5882), .n5881(n5881), .\REG.mem_8_27 (\REG.mem_8_27 ), 
            .n5880(n5880), .\REG.mem_8_26 (\REG.mem_8_26 ), .n5879(n5879), 
            .\REG.mem_8_25 (\REG.mem_8_25 ), .n5878(n5878), .n5877(n5877), 
            .n5876(n5876), .n5875(n5875), .n5874(n5874), .\REG.mem_8_20 (\REG.mem_8_20 ), 
            .n5873(n5873), .n5872(n5872), .\REG.mem_8_18 (\REG.mem_8_18 ), 
            .n5871(n5871), .n5870(n5870), .\REG.mem_8_16 (\REG.mem_8_16 ), 
            .n5869(n5869), .n5868(n5868), .\REG.mem_8_14 (\REG.mem_8_14 ), 
            .n5867(n5867), .n5866(n5866), .\REG.mem_8_12 (\REG.mem_8_12 ), 
            .n5865(n5865), .n5864(n5864), .\REG.mem_8_10 (\REG.mem_8_10 ), 
            .n5863(n5863), .\REG.mem_8_9 (\REG.mem_8_9 ), .n5862(n5862), 
            .n5861(n5861), .\REG.mem_8_7 (\REG.mem_8_7 ), .n5860(n5860), 
            .n5859(n5859), .n5858(n5858), .n5857(n5857), .\REG.mem_8_3 (\REG.mem_8_3 ), 
            .n5856(n5856), .n5855(n5855), .\REG.mem_8_1 (\REG.mem_8_1 ), 
            .n5854(n5854), .\REG.mem_8_0 (\REG.mem_8_0 ), .n5853(n5853), 
            .n5852(n5852), .n5851(n5851), .\REG.mem_7_29 (\REG.mem_7_29 ), 
            .n5850(n5850), .n5849(n5849), .n5848(n5848), .\REG.mem_7_26 (\REG.mem_7_26 ), 
            .n5847(n5847), .\REG.mem_7_25 (\REG.mem_7_25 ), .n5846(n5846), 
            .n5845(n5845), .n5844(n5844), .n5843(n5843), .n5842(n5842), 
            .\REG.mem_7_20 (\REG.mem_7_20 ), .n5841(n5841), .n5840(n5840), 
            .n5839(n5839), .n5838(n5838), .n5837(n5837), .\REG.mem_7_15 (\REG.mem_7_15 ), 
            .n5836(n5836), .\REG.mem_7_14 (\REG.mem_7_14 ), .n5835(n5835), 
            .n5834(n5834), .\REG.mem_7_12 (\REG.mem_7_12 ), .n5833(n5833), 
            .\REG.mem_7_11 (\REG.mem_7_11 ), .n5832(n5832), .n5831(n5831), 
            .n5830(n5830), .\REG.mem_7_8 (\REG.mem_7_8 ), .n5829(n5829), 
            .n5828(n5828), .n5827(n5827), .\REG.mem_7_5 (\REG.mem_7_5 ), 
            .n5826(n5826), .n5825(n5825), .\REG.mem_7_3 (\REG.mem_7_3 ), 
            .n5824(n5824), .n5823(n5823), .n5822(n5822), .n5821(n5821), 
            .n5820(n5820), .n5819(n5819), .\REG.mem_6_29 (\REG.mem_6_29 ), 
            .n5818(n5818), .n5817(n5817), .n5816(n5816), .\REG.mem_6_26 (\REG.mem_6_26 ), 
            .n5815(n5815), .\REG.mem_6_25 (\REG.mem_6_25 ), .n5814(n5814), 
            .n5813(n5813), .n5812(n5812), .n5811(n5811), .n5810(n5810), 
            .\REG.mem_6_20 (\REG.mem_6_20 ), .n5809(n5809), .n5808(n5808), 
            .n5807(n5807), .n5806(n5806), .n5805(n5805), .\REG.mem_6_15 (\REG.mem_6_15 ), 
            .n5804(n5804), .\REG.mem_6_14 (\REG.mem_6_14 ), .n5803(n5803), 
            .n5802(n5802), .\REG.mem_6_12 (\REG.mem_6_12 ), .n5801(n5801), 
            .\REG.mem_6_11 (\REG.mem_6_11 ), .n5800(n5800), .n5799(n5799), 
            .n5798(n5798), .\REG.mem_6_8 (\REG.mem_6_8 ), .n5797(n5797), 
            .n5796(n5796), .n5795(n5795), .\REG.mem_6_5 (\REG.mem_6_5 ), 
            .n5794(n5794), .n5793(n5793), .\REG.mem_6_3 (\REG.mem_6_3 ), 
            .n5792(n5792), .n5791(n5791), .n5790(n5790), .n5789(n5789), 
            .n5788(n5788), .n5600(n5600), .\REG.mem_1_3 (\REG.mem_1_3 ), 
            .n5787(n5787), .\REG.mem_5_29 (\REG.mem_5_29 ), .n25_adj_8(n25), 
            .n9(n9), .n5786(n5786), .n5785(n5785), .n5784(n5784), .\REG.mem_5_26 (\REG.mem_5_26 ), 
            .n5783(n5783), .\REG.mem_5_25 (\REG.mem_5_25 ), .n5782(n5782), 
            .\REG.mem_1_16 (\REG.mem_1_16 ), .n5781(n5781), .n5780(n5780), 
            .n5779(n5779), .n5778(n5778), .\REG.mem_5_20 (\REG.mem_5_20 ), 
            .n5777(n5777), .n5776(n5776), .n5775(n5775), .n5774(n5774), 
            .n5773(n5773), .\REG.mem_5_15 (\REG.mem_5_15 ), .n5772(n5772), 
            .\REG.mem_5_14 (\REG.mem_5_14 ), .n5771(n5771), .n5770(n5770), 
            .\REG.mem_5_12 (\REG.mem_5_12 ), .n5769(n5769), .\REG.mem_5_11 (\REG.mem_5_11 ), 
            .\REG.mem_1_25 (\REG.mem_1_25 ), .n5768(n5768), .n5767(n5767), 
            .n5766(n5766), .\REG.mem_5_8 (\REG.mem_5_8 ), .n5765(n5765), 
            .n10(n10), .n26(n26), .n5596(n5596), .n5764(n5764), .n5595(n5595), 
            .\REG.mem_1_5 (\REG.mem_1_5 ), .n5594(n5594), .n5593(n5593), 
            .n5590(n5590), .n5589(n5589), .n5588(n5588), .n5587(n5587), 
            .n5763(n5763), .\REG.mem_5_5 (\REG.mem_5_5 ), .\REG.mem_4_26 (\REG.mem_4_26 ), 
            .n5762(n5762), .n5761(n5761), .\REG.mem_5_3 (\REG.mem_5_3 ), 
            .n5760(n5760), .n5759(n5759), .n5586(n5586), .n5758(n5758), 
            .n5757(n5757), .n5756(n5756), .n5755(n5755), .\REG.mem_4_29 (\REG.mem_4_29 ), 
            .\wr_addr_nxt_c[4] (wr_addr_nxt_c[4]), .n5754(n5754), .n5753(n5753), 
            .n5752(n5752), .n5751(n5751), .\REG.mem_4_25 (\REG.mem_4_25 ), 
            .n5750(n5750), .n5749(n5749), .n5748(n5748), .n5747(n5747), 
            .n5585(n5585), .\REG.mem_1_29 (\REG.mem_1_29 ), .n5583(n5583), 
            .n5582(n5582), .n5581(n5581), .\REG.mem_1_8 (\REG.mem_1_8 ), 
            .n5580(n5580), .n5577(n5577), .n5746(n5746), .\REG.mem_4_20 (\REG.mem_4_20 ), 
            .n5745(n5745), .n5744(n5744), .n5743(n5743), .n5742(n5742), 
            .n5741(n5741), .\REG.mem_4_15 (\REG.mem_4_15 ), .n5740(n5740), 
            .\REG.mem_4_14 (\REG.mem_4_14 ), .n5739(n5739), .n5738(n5738), 
            .\REG.mem_4_12 (\REG.mem_4_12 ), .n5574(n5574), .n5572(n5572), 
            .n5571(n5571), .\REG.mem_1_11 (\REG.mem_1_11 ), .n5737(n5737), 
            .\REG.mem_4_11 (\REG.mem_4_11 ), .n5736(n5736), .n5735(n5735), 
            .n5734(n5734), .\REG.mem_4_8 (\REG.mem_4_8 ), .n5733(n5733), 
            .n5732(n5732), .n5731(n5731), .\REG.mem_4_5 (\REG.mem_4_5 ), 
            .n5730(n5730), .n5729(n5729), .\REG.mem_4_3 (\REG.mem_4_3 ), 
            .n5567(n5567), .n5565(n5565), .\REG.mem_1_20 (\REG.mem_1_20 ), 
            .n5564(n5564), .\REG.mem_1_12 (\REG.mem_1_12 ), .n5560(n5560), 
            .n5559(n5559), .\REG.mem_1_14 (\REG.mem_1_14 ), .n5558(n5558), 
            .\REG.mem_1_15 (\REG.mem_1_15 ), .n5557(n5557), .n5556(n5556), 
            .n5555(n5555), .n5554(n5554), .n5551(n5551), .n5550(n5550), 
            .n5728(n5728), .n5727(n5727), .n5726(n5726), .n11(n11), 
            .n27(n27)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(579[21] 595[2])
    SB_LUT4 i1937_2_lut_3_lut_4_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(reset_all_w), .I3(wr_addr_r_adj_1517[0]), .O(n8_adj_1418));
    defparam i1937_2_lut_3_lut_4_lut.LUT_INIT = 16'h0df2;
    SB_LUT4 i4507_3_lut (.I0(\REG.mem_11_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n22), .I3(GND_net), .O(n5981));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4506_3_lut (.I0(\REG.mem_11_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n22), .I3(GND_net), .O(n5980));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4505_3_lut (.I0(\REG.mem_11_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n22), .I3(GND_net), .O(n5979));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4504_3_lut (.I0(\REG.mem_11_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n22), .I3(GND_net), .O(n5978));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4503_3_lut (.I0(\REG.mem_11_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n22), .I3(GND_net), .O(n5977));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4502_3_lut (.I0(\REG.mem_11_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n22), .I3(GND_net), .O(n5976));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4501_3_lut (.I0(\REG.mem_11_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n22), .I3(GND_net), .O(n5975));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4500_3_lut (.I0(\REG.mem_11_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n22), .I3(GND_net), .O(n5974));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4499_3_lut (.I0(\REG.mem_11_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n22), .I3(GND_net), .O(n5973));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4498_3_lut (.I0(\REG.mem_11_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n22), .I3(GND_net), .O(n5972));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4497_3_lut (.I0(\REG.mem_11_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n22), .I3(GND_net), .O(n5971));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4496_3_lut (.I0(\REG.mem_11_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n22), .I3(GND_net), .O(n5970));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4141_3_lut (.I0(tx_addr_byte[0]), .I1(tx_data_byte[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5615));   // src/top.v(1165[8] 1232[4])
    defparam i4141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4495_3_lut (.I0(\REG.mem_11_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n22), .I3(GND_net), .O(n5969));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4494_3_lut (.I0(\REG.mem_11_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n22), .I3(GND_net), .O(n5968));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4493_3_lut (.I0(\REG.mem_11_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n22), .I3(GND_net), .O(n5967));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4493_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4492_3_lut (.I0(\REG.mem_11_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n22), .I3(GND_net), .O(n5966));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4491_3_lut (.I0(\REG.mem_11_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n22), .I3(GND_net), .O(n5965));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4490_3_lut (.I0(\REG.mem_11_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n22), .I3(GND_net), .O(n5964));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4489_3_lut (.I0(\REG.mem_11_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n22), .I3(GND_net), .O(n5963));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4488_3_lut (.I0(\REG.mem_11_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n22), .I3(GND_net), .O(n5962));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4487_3_lut (.I0(\REG.mem_11_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n22), .I3(GND_net), .O(n5961));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4486_3_lut (.I0(\REG.mem_11_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n22), .I3(GND_net), .O(n5960));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4485_3_lut (.I0(\REG.mem_11_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n22), .I3(GND_net), .O(n5959));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4484_3_lut (.I0(\REG.mem_11_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n22), .I3(GND_net), .O(n5958));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4484_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4483_3_lut (.I0(\REG.mem_11_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n22), .I3(GND_net), .O(n5957));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4482_3_lut (.I0(\REG.mem_11_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n22), .I3(GND_net), .O(n5956));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4481_3_lut (.I0(\REG.mem_11_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n22), .I3(GND_net), .O(n5955));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4480_3_lut (.I0(\REG.mem_11_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n22), .I3(GND_net), .O(n5954));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4479_3_lut (.I0(\REG.mem_11_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n22), .I3(GND_net), .O(n5953));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_125 (.I0(buffer_switch_done_latched), .I1(n1013), 
            .I2(n934), .I3(GND_net), .O(n12261));
    defparam i1_3_lut_adj_125.LUT_INIT = 16'heaea;
    SB_LUT4 i4478_3_lut (.I0(\REG.mem_11_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n22), .I3(GND_net), .O(n5952));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4477_3_lut (.I0(\REG.mem_11_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n22), .I3(GND_net), .O(n5951));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4476_3_lut (.I0(\REG.mem_11_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n22), .I3(GND_net), .O(n5950));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4475_3_lut (.I0(\REG.mem_10_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n23), .I3(GND_net), .O(n5949));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4474_3_lut (.I0(\REG.mem_10_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n23), .I3(GND_net), .O(n5948));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4473_3_lut (.I0(\REG.mem_10_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n23), .I3(GND_net), .O(n5947));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4472_3_lut (.I0(\REG.mem_10_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n23), .I3(GND_net), .O(n5946));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4471_3_lut (.I0(\REG.mem_10_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n23), .I3(GND_net), .O(n5945));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4470_3_lut (.I0(\REG.mem_10_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n23), .I3(GND_net), .O(n5944));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4469_3_lut (.I0(\REG.mem_10_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n23), .I3(GND_net), .O(n5943));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4468_3_lut (.I0(\REG.mem_10_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n23), .I3(GND_net), .O(n5942));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4137_3_lut (.I0(\REG.mem_1_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n32), .I3(GND_net), .O(n5611));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4136_3_lut (.I0(\REG.mem_1_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n32), .I3(GND_net), .O(n5610));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4467_3_lut (.I0(\REG.mem_10_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n23), .I3(GND_net), .O(n5941));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4466_3_lut (.I0(\REG.mem_10_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n23), .I3(GND_net), .O(n5940));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4466_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4465_3_lut (.I0(\REG.mem_10_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n23), .I3(GND_net), .O(n5939));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4464_3_lut (.I0(\REG.mem_10_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n23), .I3(GND_net), .O(n5938));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4463_3_lut (.I0(\REG.mem_10_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n23), .I3(GND_net), .O(n5937));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_126 (.I0(reset_all_w), .I1(n12964), .I2(n24_adj_1443), 
            .I3(n4_adj_1441), .O(n12836));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_adj_126.LUT_INIT = 16'hfbfa;
    SB_LUT4 i10857_4_lut (.I0(rd_addr_p1_w_adj_1522[2]), .I1(rd_addr_p1_w_adj_1522[1]), 
            .I2(wr_addr_r_adj_1517[2]), .I3(wr_addr_r_adj_1517[1]), .O(n12964));
    defparam i10857_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_3_lut_adj_127 (.I0(is_fifo_empty_flag), .I1(fifo_write_cmd), 
            .I2(n32_adj_1440), .I3(GND_net), .O(n24_adj_1443));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_3_lut_adj_127.LUT_INIT = 16'h2020;
    SB_LUT4 i1_4_lut_adj_128 (.I0(rd_addr_r_adj_1520[1]), .I1(rd_addr_r_adj_1520[0]), 
            .I2(wr_addr_r_adj_1517[1]), .I3(wr_addr_r_adj_1517[0]), .O(n32_adj_1440));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_adj_128.LUT_INIT = 16'h8421;
    SB_LUT4 i4134_3_lut (.I0(\REG.mem_1_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n32), .I3(GND_net), .O(n5608));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4130_3_lut (.I0(\REG.mem_1_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n32), .I3(GND_net), .O(n5604));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4129_3_lut (.I0(\REG.mem_1_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n32), .I3(GND_net), .O(n5603));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4128_3_lut (.I0(\REG.mem_1_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n32), .I3(GND_net), .O(n5602));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4462_3_lut (.I0(\REG.mem_10_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n23), .I3(GND_net), .O(n5936));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4461_3_lut (.I0(\REG.mem_10_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n23), .I3(GND_net), .O(n5935));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4460_3_lut (.I0(\REG.mem_10_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n23), .I3(GND_net), .O(n5934));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4459_3_lut (.I0(\REG.mem_10_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n23), .I3(GND_net), .O(n5933));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4458_3_lut (.I0(\REG.mem_10_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n23), .I3(GND_net), .O(n5932));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4457_3_lut (.I0(\REG.mem_10_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n23), .I3(GND_net), .O(n5931));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4456_3_lut (.I0(\REG.mem_10_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n23), .I3(GND_net), .O(n5930));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4455_3_lut (.I0(\REG.mem_10_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n23), .I3(GND_net), .O(n5929));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4454_3_lut (.I0(\REG.mem_10_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n23), .I3(GND_net), .O(n5928));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4453_3_lut (.I0(\REG.mem_10_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n23), .I3(GND_net), .O(n5927));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4452_3_lut (.I0(\REG.mem_10_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n23), .I3(GND_net), .O(n5926));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4451_3_lut (.I0(\REG.mem_10_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n23), .I3(GND_net), .O(n5925));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4450_3_lut (.I0(\REG.mem_10_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n23), .I3(GND_net), .O(n5924));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4449_3_lut (.I0(\REG.mem_10_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n23), .I3(GND_net), .O(n5923));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4448_3_lut (.I0(\REG.mem_10_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n23), .I3(GND_net), .O(n5922));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4447_3_lut (.I0(\REG.mem_10_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n23), .I3(GND_net), .O(n5921));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4446_3_lut (.I0(\REG.mem_10_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n23), .I3(GND_net), .O(n5920));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4445_3_lut (.I0(\REG.mem_10_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n23), .I3(GND_net), .O(n5919));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4444_3_lut (.I0(\REG.mem_10_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n23), .I3(GND_net), .O(n5918));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4443_3_lut (.I0(\REG.mem_9_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n24), .I3(GND_net), .O(n5917));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4442_3_lut (.I0(\REG.mem_9_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n24), .I3(GND_net), .O(n5916));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4441_3_lut (.I0(\REG.mem_9_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n24), .I3(GND_net), .O(n5915));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4440_3_lut (.I0(\REG.mem_9_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n24), .I3(GND_net), .O(n5914));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4439_3_lut (.I0(\REG.mem_9_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n24), .I3(GND_net), .O(n5913));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4438_3_lut (.I0(\REG.mem_9_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n24), .I3(GND_net), .O(n5912));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4437_3_lut (.I0(\REG.mem_9_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n24), .I3(GND_net), .O(n5911));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4436_3_lut (.I0(\REG.mem_9_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n24), .I3(GND_net), .O(n5910));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4435_3_lut (.I0(\REG.mem_9_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n24), .I3(GND_net), .O(n5909));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4434_3_lut (.I0(\REG.mem_9_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n24), .I3(GND_net), .O(n5908));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4433_3_lut (.I0(\REG.mem_9_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n24), .I3(GND_net), .O(n5907));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4432_3_lut (.I0(\REG.mem_9_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n24), .I3(GND_net), .O(n5906));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4431_3_lut (.I0(\REG.mem_9_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n24), .I3(GND_net), .O(n5905));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4430_3_lut (.I0(\REG.mem_9_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n24), .I3(GND_net), .O(n5904));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4429_3_lut (.I0(\REG.mem_9_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n24), .I3(GND_net), .O(n5903));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4429_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4428_3_lut (.I0(\REG.mem_9_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n24), .I3(GND_net), .O(n5902));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4427_3_lut (.I0(\REG.mem_9_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n24), .I3(GND_net), .O(n5901));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4426_3_lut (.I0(\REG.mem_9_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n24), .I3(GND_net), .O(n5900));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4425_3_lut (.I0(\REG.mem_9_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n24), .I3(GND_net), .O(n5899));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4424_3_lut (.I0(\REG.mem_9_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n24), .I3(GND_net), .O(n5898));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4423_3_lut (.I0(\REG.mem_9_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n24), .I3(GND_net), .O(n5897));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4422_3_lut (.I0(\REG.mem_9_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n24), .I3(GND_net), .O(n5896));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4421_3_lut (.I0(\REG.mem_9_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n24), .I3(GND_net), .O(n5895));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4420_3_lut (.I0(\REG.mem_9_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n24), .I3(GND_net), .O(n5894));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4419_3_lut (.I0(\REG.mem_9_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n24), .I3(GND_net), .O(n5893));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4418_3_lut (.I0(\REG.mem_9_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n24), .I3(GND_net), .O(n5892));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4417_3_lut (.I0(\REG.mem_9_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n24), .I3(GND_net), .O(n5891));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4416_3_lut (.I0(\REG.mem_9_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n24), .I3(GND_net), .O(n5890));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4415_3_lut (.I0(\REG.mem_9_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n24), .I3(GND_net), .O(n5889));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4414_3_lut (.I0(\REG.mem_9_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n24), .I3(GND_net), .O(n5888));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4413_3_lut (.I0(\REG.mem_9_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n24), .I3(GND_net), .O(n5887));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4412_3_lut (.I0(\REG.mem_9_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n24), .I3(GND_net), .O(n5886));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4411_3_lut (.I0(\REG.mem_8_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n25), .I3(GND_net), .O(n5885));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4410_3_lut (.I0(\REG.mem_8_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n25), .I3(GND_net), .O(n5884));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4409_3_lut (.I0(\REG.mem_8_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n25), .I3(GND_net), .O(n5883));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4408_3_lut (.I0(\REG.mem_8_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n25), .I3(GND_net), .O(n5882));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4407_3_lut (.I0(\REG.mem_8_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n25), .I3(GND_net), .O(n5881));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4406_3_lut (.I0(\REG.mem_8_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n25), .I3(GND_net), .O(n5880));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4405_3_lut (.I0(\REG.mem_8_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n25), .I3(GND_net), .O(n5879));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4404_3_lut (.I0(\REG.mem_8_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n25), .I3(GND_net), .O(n5878));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4404_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4403_3_lut (.I0(\REG.mem_8_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n25), .I3(GND_net), .O(n5877));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4402_3_lut (.I0(\REG.mem_8_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n25), .I3(GND_net), .O(n5876));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4401_3_lut (.I0(\REG.mem_8_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n25), .I3(GND_net), .O(n5875));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4400_3_lut (.I0(\REG.mem_8_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n25), .I3(GND_net), .O(n5874));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4399_3_lut (.I0(\REG.mem_8_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n25), .I3(GND_net), .O(n5873));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4398_3_lut (.I0(\REG.mem_8_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n25), .I3(GND_net), .O(n5872));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4397_3_lut (.I0(\REG.mem_8_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n25), .I3(GND_net), .O(n5871));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4396_3_lut (.I0(\REG.mem_8_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n25), .I3(GND_net), .O(n5870));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4395_3_lut (.I0(\REG.mem_8_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n25), .I3(GND_net), .O(n5869));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4394_3_lut (.I0(\REG.mem_8_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n25), .I3(GND_net), .O(n5868));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4393_3_lut (.I0(\REG.mem_8_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n25), .I3(GND_net), .O(n5867));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4392_3_lut (.I0(\REG.mem_8_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n25), .I3(GND_net), .O(n5866));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4391_3_lut (.I0(\REG.mem_8_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n25), .I3(GND_net), .O(n5865));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4390_3_lut (.I0(\REG.mem_8_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n25), .I3(GND_net), .O(n5864));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4389_3_lut (.I0(\REG.mem_8_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n25), .I3(GND_net), .O(n5863));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4388_3_lut (.I0(\REG.mem_8_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n25), .I3(GND_net), .O(n5862));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4387_3_lut (.I0(\REG.mem_8_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n25), .I3(GND_net), .O(n5861));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4386_3_lut (.I0(\REG.mem_8_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n25), .I3(GND_net), .O(n5860));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4385_3_lut (.I0(\REG.mem_8_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n25), .I3(GND_net), .O(n5859));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4384_3_lut (.I0(\REG.mem_8_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n25), .I3(GND_net), .O(n5858));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4383_3_lut (.I0(\REG.mem_8_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n25), .I3(GND_net), .O(n5857));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4382_3_lut (.I0(\REG.mem_8_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n25), .I3(GND_net), .O(n5856));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4381_3_lut (.I0(\REG.mem_8_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n25), .I3(GND_net), .O(n5855));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4380_3_lut (.I0(\REG.mem_8_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n25), .I3(GND_net), .O(n5854));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4379_3_lut (.I0(\REG.mem_7_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n26), .I3(GND_net), .O(n5853));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4378_3_lut (.I0(\REG.mem_7_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n26), .I3(GND_net), .O(n5852));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4377_3_lut (.I0(\REG.mem_7_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n26), .I3(GND_net), .O(n5851));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4376_3_lut (.I0(\REG.mem_7_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n26), .I3(GND_net), .O(n5850));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4375_3_lut (.I0(\REG.mem_7_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n26), .I3(GND_net), .O(n5849));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4374_3_lut (.I0(\REG.mem_7_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n26), .I3(GND_net), .O(n5848));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4373_3_lut (.I0(\REG.mem_7_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n26), .I3(GND_net), .O(n5847));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4372_3_lut (.I0(\REG.mem_7_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n26), .I3(GND_net), .O(n5846));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4371_3_lut (.I0(\REG.mem_7_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n26), .I3(GND_net), .O(n5845));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4370_3_lut (.I0(\REG.mem_7_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n26), .I3(GND_net), .O(n5844));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4369_3_lut (.I0(\REG.mem_7_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n26), .I3(GND_net), .O(n5843));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4368_3_lut (.I0(\REG.mem_7_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n26), .I3(GND_net), .O(n5842));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4367_3_lut (.I0(\REG.mem_7_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n26), .I3(GND_net), .O(n5841));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4366_3_lut (.I0(\REG.mem_7_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n26), .I3(GND_net), .O(n5840));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4365_3_lut (.I0(\REG.mem_7_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n26), .I3(GND_net), .O(n5839));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4364_3_lut (.I0(\REG.mem_7_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n26), .I3(GND_net), .O(n5838));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4363_3_lut (.I0(\REG.mem_7_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n26), .I3(GND_net), .O(n5837));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4362_3_lut (.I0(\REG.mem_7_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n26), .I3(GND_net), .O(n5836));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4361_3_lut (.I0(\REG.mem_7_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n26), .I3(GND_net), .O(n5835));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4360_3_lut (.I0(\REG.mem_7_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n26), .I3(GND_net), .O(n5834));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4359_3_lut (.I0(\REG.mem_7_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n26), .I3(GND_net), .O(n5833));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4358_3_lut (.I0(\REG.mem_7_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n26), .I3(GND_net), .O(n5832));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4357_3_lut (.I0(\REG.mem_7_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n26), .I3(GND_net), .O(n5831));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4356_3_lut (.I0(\REG.mem_7_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n26), .I3(GND_net), .O(n5830));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4355_3_lut (.I0(\REG.mem_7_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n26), .I3(GND_net), .O(n5829));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4354_3_lut (.I0(\REG.mem_7_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n26), .I3(GND_net), .O(n5828));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4353_3_lut (.I0(\REG.mem_7_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n26), .I3(GND_net), .O(n5827));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4352_3_lut (.I0(\REG.mem_7_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n26), .I3(GND_net), .O(n5826));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4351_3_lut (.I0(\REG.mem_7_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n26), .I3(GND_net), .O(n5825));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4350_3_lut (.I0(\REG.mem_7_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n26), .I3(GND_net), .O(n5824));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4349_3_lut (.I0(\REG.mem_7_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n26), .I3(GND_net), .O(n5823));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4348_3_lut (.I0(\REG.mem_7_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n26), .I3(GND_net), .O(n5822));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4347_3_lut (.I0(\REG.mem_6_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n27), .I3(GND_net), .O(n5821));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4346_3_lut (.I0(\REG.mem_6_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n27), .I3(GND_net), .O(n5820));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4345_3_lut (.I0(\REG.mem_6_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n27), .I3(GND_net), .O(n5819));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4344_3_lut (.I0(\REG.mem_6_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n27), .I3(GND_net), .O(n5818));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4343_3_lut (.I0(\REG.mem_6_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n27), .I3(GND_net), .O(n5817));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4342_3_lut (.I0(\REG.mem_6_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n27), .I3(GND_net), .O(n5816));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4341_3_lut (.I0(\REG.mem_6_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n27), .I3(GND_net), .O(n5815));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4340_3_lut (.I0(\REG.mem_6_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n27), .I3(GND_net), .O(n5814));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4339_3_lut (.I0(\REG.mem_6_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n27), .I3(GND_net), .O(n5813));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4338_3_lut (.I0(\REG.mem_6_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n27), .I3(GND_net), .O(n5812));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4337_3_lut (.I0(\REG.mem_6_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n27), .I3(GND_net), .O(n5811));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4336_3_lut (.I0(\REG.mem_6_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n27), .I3(GND_net), .O(n5810));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4335_3_lut (.I0(\REG.mem_6_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n27), .I3(GND_net), .O(n5809));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4334_3_lut (.I0(\REG.mem_6_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n27), .I3(GND_net), .O(n5808));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4333_3_lut (.I0(\REG.mem_6_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n27), .I3(GND_net), .O(n5807));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4332_3_lut (.I0(\REG.mem_6_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n27), .I3(GND_net), .O(n5806));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4331_3_lut (.I0(\REG.mem_6_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n27), .I3(GND_net), .O(n5805));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4330_3_lut (.I0(\REG.mem_6_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n27), .I3(GND_net), .O(n5804));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4329_3_lut (.I0(\REG.mem_6_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n27), .I3(GND_net), .O(n5803));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4328_3_lut (.I0(\REG.mem_6_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n27), .I3(GND_net), .O(n5802));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4327_3_lut (.I0(\REG.mem_6_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n27), .I3(GND_net), .O(n5801));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4326_3_lut (.I0(\REG.mem_6_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n27), .I3(GND_net), .O(n5800));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4325_3_lut (.I0(\REG.mem_6_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n27), .I3(GND_net), .O(n5799));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4324_3_lut (.I0(\REG.mem_6_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n27), .I3(GND_net), .O(n5798));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4323_3_lut (.I0(\REG.mem_6_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n27), .I3(GND_net), .O(n5797));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4322_3_lut (.I0(\REG.mem_6_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n27), .I3(GND_net), .O(n5796));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4321_3_lut (.I0(\REG.mem_6_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n27), .I3(GND_net), .O(n5795));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4320_3_lut (.I0(\REG.mem_6_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n27), .I3(GND_net), .O(n5794));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4319_3_lut (.I0(\REG.mem_6_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n27), .I3(GND_net), .O(n5793));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4318_3_lut (.I0(\REG.mem_6_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n27), .I3(GND_net), .O(n5792));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4317_3_lut (.I0(\REG.mem_6_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n27), .I3(GND_net), .O(n5791));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4316_3_lut (.I0(\REG.mem_6_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n27), .I3(GND_net), .O(n5790));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4315_3_lut (.I0(\REG.mem_5_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n28), .I3(GND_net), .O(n5789));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4314_3_lut (.I0(\REG.mem_5_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n28), .I3(GND_net), .O(n5788));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4126_3_lut (.I0(\REG.mem_1_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n32), .I3(GND_net), .O(n5600));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4313_3_lut (.I0(\REG.mem_5_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n28), .I3(GND_net), .O(n5787));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4312_3_lut (.I0(\REG.mem_5_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n28), .I3(GND_net), .O(n5786));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4311_3_lut (.I0(\REG.mem_5_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n28), .I3(GND_net), .O(n5785));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4310_3_lut (.I0(\REG.mem_5_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n28), .I3(GND_net), .O(n5784));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4309_3_lut (.I0(\REG.mem_5_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n28), .I3(GND_net), .O(n5783));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4308_3_lut (.I0(\REG.mem_5_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n28), .I3(GND_net), .O(n5782));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4307_3_lut (.I0(\REG.mem_5_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n28), .I3(GND_net), .O(n5781));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4306_3_lut (.I0(\REG.mem_5_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n28), .I3(GND_net), .O(n5780));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4305_3_lut (.I0(\REG.mem_5_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n28), .I3(GND_net), .O(n5779));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4304_3_lut (.I0(\REG.mem_5_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n28), .I3(GND_net), .O(n5778));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4303_3_lut (.I0(\REG.mem_5_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n28), .I3(GND_net), .O(n5777));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4302_3_lut (.I0(\REG.mem_5_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n28), .I3(GND_net), .O(n5776));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4301_3_lut (.I0(\REG.mem_5_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n28), .I3(GND_net), .O(n5775));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4300_3_lut (.I0(\REG.mem_5_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n28), .I3(GND_net), .O(n5774));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4299_3_lut (.I0(\REG.mem_5_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n28), .I3(GND_net), .O(n5773));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4298_3_lut (.I0(\REG.mem_5_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n28), .I3(GND_net), .O(n5772));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4297_3_lut (.I0(\REG.mem_5_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n28), .I3(GND_net), .O(n5771));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4296_3_lut (.I0(\REG.mem_5_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n28), .I3(GND_net), .O(n5770));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4295_3_lut (.I0(\REG.mem_5_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n28), .I3(GND_net), .O(n5769));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4294_3_lut (.I0(\REG.mem_5_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n28), .I3(GND_net), .O(n5768));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4293_3_lut (.I0(\REG.mem_5_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n28), .I3(GND_net), .O(n5767));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4292_3_lut (.I0(\REG.mem_5_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n28), .I3(GND_net), .O(n5766));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4291_3_lut (.I0(\REG.mem_5_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n28), .I3(GND_net), .O(n5765));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4122_3_lut (.I0(\REG.mem_1_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n32), .I3(GND_net), .O(n5596));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4290_3_lut (.I0(\REG.mem_5_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n28), .I3(GND_net), .O(n5764));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4121_3_lut (.I0(\REG.mem_1_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n32), .I3(GND_net), .O(n5595));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4120_3_lut (.I0(\REG.mem_1_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n32), .I3(GND_net), .O(n5594));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4119_3_lut (.I0(\REG.mem_1_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n32), .I3(GND_net), .O(n5593));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4118_2_lut (.I0(uart_rx_complete_prev), .I1(debug_led3), .I2(GND_net), 
            .I3(GND_net), .O(n5592));   // src/top.v(1156[8] 1162[4])
    defparam i4118_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4116_3_lut (.I0(\REG.mem_1_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n32), .I3(GND_net), .O(n5590));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4115_3_lut (.I0(\REG.mem_1_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n32), .I3(GND_net), .O(n5589));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4114_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5588));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4114_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4113_3_lut (.I0(\REG.mem_1_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n32), .I3(GND_net), .O(n5587));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4289_3_lut (.I0(\REG.mem_5_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n28), .I3(GND_net), .O(n5763));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4288_3_lut (.I0(\REG.mem_5_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n28), .I3(GND_net), .O(n5762));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4287_3_lut (.I0(\REG.mem_5_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n28), .I3(GND_net), .O(n5761));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4286_3_lut (.I0(\REG.mem_5_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n28), .I3(GND_net), .O(n5760));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4285_3_lut (.I0(\REG.mem_5_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n28), .I3(GND_net), .O(n5759));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4112_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5586));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4112_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4284_3_lut (.I0(\REG.mem_5_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n28), .I3(GND_net), .O(n5758));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4283_3_lut (.I0(\REG.mem_4_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n29), .I3(GND_net), .O(n5757));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4282_3_lut (.I0(\REG.mem_4_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n29), .I3(GND_net), .O(n5756));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_129 (.I0(reset_clk_counter[3]), .I1(reset_clk_counter[2]), 
            .I2(n12040), .I3(GND_net), .O(n12308));
    defparam i1_3_lut_adj_129.LUT_INIT = 16'ha9a9;
    SB_LUT4 i4281_3_lut (.I0(\REG.mem_4_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n29), .I3(GND_net), .O(n5755));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4280_3_lut (.I0(\REG.mem_4_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n29), .I3(GND_net), .O(n5754));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4279_3_lut (.I0(\REG.mem_4_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n29), .I3(GND_net), .O(n5753));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4278_3_lut (.I0(\REG.mem_4_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n29), .I3(GND_net), .O(n5752));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4277_3_lut (.I0(\REG.mem_4_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n29), .I3(GND_net), .O(n5751));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4276_3_lut (.I0(\REG.mem_4_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n29), .I3(GND_net), .O(n5750));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4275_3_lut (.I0(\REG.mem_4_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n29), .I3(GND_net), .O(n5749));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4274_3_lut (.I0(\REG.mem_4_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n29), .I3(GND_net), .O(n5748));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4274_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4273_3_lut (.I0(\REG.mem_4_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n29), .I3(GND_net), .O(n5747));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4111_3_lut (.I0(\REG.mem_1_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n32), .I3(GND_net), .O(n5585));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4109_3_lut (.I0(\REG.mem_1_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n32), .I3(GND_net), .O(n5583));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4108_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5582));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4108_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4107_3_lut (.I0(\REG.mem_1_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n32), .I3(GND_net), .O(n5581));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4106_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5580));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4106_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4104_3_lut (.I0(rx_buf_byte[0]), .I1(rx_shift_reg[0]), .I2(n3963), 
            .I3(GND_net), .O(n5578));   // src/spi.v(76[8] 221[4])
    defparam i4104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4103_3_lut (.I0(\REG.mem_1_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n32), .I3(GND_net), .O(n5577));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4272_3_lut (.I0(\REG.mem_4_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n29), .I3(GND_net), .O(n5746));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4271_3_lut (.I0(\REG.mem_4_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n29), .I3(GND_net), .O(n5745));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4270_3_lut (.I0(\REG.mem_4_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n29), .I3(GND_net), .O(n5744));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4269_3_lut (.I0(\REG.mem_4_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n29), .I3(GND_net), .O(n5743));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4268_3_lut (.I0(\REG.mem_4_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n29), .I3(GND_net), .O(n5742));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4267_3_lut (.I0(\REG.mem_4_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n29), .I3(GND_net), .O(n5741));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4266_3_lut (.I0(\REG.mem_4_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n29), .I3(GND_net), .O(n5740));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4265_3_lut (.I0(\REG.mem_4_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n29), .I3(GND_net), .O(n5739));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4264_3_lut (.I0(\REG.mem_4_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n29), .I3(GND_net), .O(n5738));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4102_3_lut (.I0(r_Tx_Data[0]), .I1(fifo_temp_output[0]), .I2(n4314), 
            .I3(GND_net), .O(n5576));   // src/uart_tx.v(38[10] 141[8])
    defparam i4102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4100_3_lut (.I0(\REG.mem_1_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n32), .I3(GND_net), .O(n5574));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4099_2_lut (.I0(bluejay_data_out_31__N_920), .I1(bluejay_data_out_31__N_921), 
            .I2(GND_net), .I3(GND_net), .O(n5573));   // src/bluejay_data.v(134[8] 156[4])
    defparam i4099_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4098_3_lut (.I0(\REG.mem_1_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n32), .I3(GND_net), .O(n5572));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4097_3_lut (.I0(\REG.mem_1_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n32), .I3(GND_net), .O(n5571));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4263_3_lut (.I0(\REG.mem_4_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n29), .I3(GND_net), .O(n5737));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4262_3_lut (.I0(\REG.mem_4_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n29), .I3(GND_net), .O(n5736));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4261_3_lut (.I0(\REG.mem_4_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n29), .I3(GND_net), .O(n5735));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4260_3_lut (.I0(\REG.mem_4_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n29), .I3(GND_net), .O(n5734));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4259_3_lut (.I0(\REG.mem_4_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n29), .I3(GND_net), .O(n5733));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4258_3_lut (.I0(\REG.mem_4_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n29), .I3(GND_net), .O(n5732));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4257_3_lut (.I0(\REG.mem_4_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n29), .I3(GND_net), .O(n5731));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4256_3_lut (.I0(\REG.mem_4_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n29), .I3(GND_net), .O(n5730));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4255_3_lut (.I0(\REG.mem_4_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n29), .I3(GND_net), .O(n5729));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4093_3_lut (.I0(\REG.mem_1_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n32), .I3(GND_net), .O(n5567));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_130 (.I0(n63), .I1(state[1]), .I2(state[3]), 
            .I3(n12882), .O(n12884));   // src/timing_controller.v(160[5] 229[12])
    defparam i3_4_lut_adj_130.LUT_INIT = 16'h0400;
    SB_LUT4 i4091_3_lut (.I0(\REG.mem_1_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n32), .I3(GND_net), .O(n5565));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4090_3_lut (.I0(\REG.mem_1_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n32), .I3(GND_net), .O(n5564));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1936_2_lut_3_lut_4_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(reset_all_w), .I3(rd_addr_r_adj_1520[0]), .O(n8));
    defparam i1936_2_lut_3_lut_4_lut.LUT_INIT = 16'h0df2;
    SB_LUT4 i4086_3_lut (.I0(\REG.mem_1_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n32), .I3(GND_net), .O(n5560));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4085_3_lut (.I0(\REG.mem_1_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n32), .I3(GND_net), .O(n5559));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4084_3_lut (.I0(\REG.mem_1_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n32), .I3(GND_net), .O(n5558));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4083_3_lut (.I0(\REG.mem_1_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n32), .I3(GND_net), .O(n5557));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4082_3_lut (.I0(\REG.mem_1_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n32), .I3(GND_net), .O(n5556));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4081_3_lut (.I0(\REG.mem_1_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n32), .I3(GND_net), .O(n5555));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4078_3_lut (.I0(tx_data_byte[0]), .I1(pc_data_rx[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5552));   // src/top.v(1165[8] 1232[4])
    defparam i4078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4077_3_lut (.I0(\REG.mem_1_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n32), .I3(GND_net), .O(n5551));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4076_3_lut (.I0(\REG.mem_1_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n32), .I3(GND_net), .O(n5550));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4254_3_lut (.I0(\REG.mem_4_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n29), .I3(GND_net), .O(n5728));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4253_3_lut (.I0(\REG.mem_4_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n29), .I3(GND_net), .O(n5727));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4252_3_lut (.I0(\REG.mem_4_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n29), .I3(GND_net), .O(n5726));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(reset_all_w), .I3(rd_fifo_en_prev_r), .O(n5086));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff2;
    FIFO_Quad_Word tx_fifo (.n8(n8), .rd_addr_r({rd_addr_r_adj_1520}), .SLM_CLK_c(SLM_CLK_c), 
            .reset_all_w(reset_all_w), .wr_addr_r({wr_addr_r_adj_1517}), 
            .rx_buf_byte({rx_buf_byte}), .n4446(n4446), .GND_net(GND_net), 
            .\wr_addr_p1_w[2] (wr_addr_p1_w_adj_1519[2]), .n12215(n12215), 
            .rd_fifo_en_w(rd_fifo_en_w), .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r [0]), 
            .n8_adj_2(n8_adj_1418), .n5599(n5599), .n5607(n5607), .n12439(n12439), 
            .VCC_net(VCC_net), .is_tx_fifo_full_flag(is_tx_fifo_full_flag), 
            .n5645(n5645), .\fifo_temp_output[7] (fifo_temp_output[7]), 
            .n5648(n5648), .\fifo_temp_output[6] (fifo_temp_output[6]), 
            .n5653(n5653), .\fifo_temp_output[5] (fifo_temp_output[5]), 
            .n6947(n6947), .\fifo_temp_output[0] (fifo_temp_output[0]), 
            .n5656(n5656), .\fifo_temp_output[4] (fifo_temp_output[4]), 
            .n5659(n5659), .\fifo_temp_output[3] (fifo_temp_output[3]), 
            .n5662(n5662), .\fifo_temp_output[2] (fifo_temp_output[2]), 
            .n5665(n5665), .\fifo_temp_output[1] (fifo_temp_output[1]), 
            .n6923(n6923), .n6920(n6920), .fifo_write_cmd(fifo_write_cmd), 
            .wr_fifo_en_w(wr_fifo_en_w_adj_1416), .n5636(n5636), .rd_fifo_en_prev_r(rd_fifo_en_prev_r), 
            .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r [1]), .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r [2]), 
            .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r [3]), .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r [4]), 
            .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r [5]), .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r [6]), 
            .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r [7]), .n12836(n12836), 
            .is_fifo_empty_flag(is_fifo_empty_flag), .fifo_read_cmd(fifo_read_cmd), 
            .\rd_addr_p1_w[2] (rd_addr_p1_w_adj_1522[2]), .\rd_addr_p1_w[1] (rd_addr_p1_w_adj_1522[1])) /* synthesis syn_module_defined=1 */ ;   // src/top.v(1024[16] 1040[2])
    SB_LUT4 i1_4_lut_4_lut (.I0(is_tx_fifo_full_flag), .I1(n12938), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h2222;
    fifo_sc_32_lut_gen fifo_sc_32_lut_gen_inst (.DEBUG_9_c_0(DEBUG_9_c_0), 
            .SLM_CLK_c(SLM_CLK_c), .\dc32_fifo_data_out[31] (dc32_fifo_data_out[31]), 
            .\dc32_fifo_data_out[30] (dc32_fifo_data_out[30]), .\dc32_fifo_data_out[29] (dc32_fifo_data_out[29]), 
            .\dc32_fifo_data_out[28] (dc32_fifo_data_out[28]), .\dc32_fifo_data_out[27] (dc32_fifo_data_out[27]), 
            .\dc32_fifo_data_out[26] (dc32_fifo_data_out[26]), .\dc32_fifo_data_out[25] (dc32_fifo_data_out[25]), 
            .\dc32_fifo_data_out[24] (dc32_fifo_data_out[24]), .\dc32_fifo_data_out[23] (dc32_fifo_data_out[23]), 
            .sc32_fifo_almost_empty(sc32_fifo_almost_empty), .reset_all(reset_all), 
            .\dc32_fifo_data_out[22] (dc32_fifo_data_out[22]), .\dc32_fifo_data_out[21] (dc32_fifo_data_out[21]), 
            .\dc32_fifo_data_out[20] (dc32_fifo_data_out[20]), .\dc32_fifo_data_out[19] (dc32_fifo_data_out[19]), 
            .\dc32_fifo_data_out[18] (dc32_fifo_data_out[18]), .\dc32_fifo_data_out[17] (dc32_fifo_data_out[17]), 
            .\dc32_fifo_data_out[16] (dc32_fifo_data_out[16]), .\dc32_fifo_data_out[15] (dc32_fifo_data_out[15]), 
            .\dc32_fifo_data_out[14] (dc32_fifo_data_out[14]), .\dc32_fifo_data_out[13] (dc32_fifo_data_out[13]), 
            .\dc32_fifo_data_out[12] (dc32_fifo_data_out[12]), .\dc32_fifo_data_out[11] (dc32_fifo_data_out[11]), 
            .\dc32_fifo_data_out[10] (dc32_fifo_data_out[10]), .\dc32_fifo_data_out[9] (dc32_fifo_data_out[9]), 
            .\dc32_fifo_data_out[8] (dc32_fifo_data_out[8]), .\dc32_fifo_data_out[7] (dc32_fifo_data_out[7]), 
            .\dc32_fifo_data_out[6] (dc32_fifo_data_out[6]), .GND_net(GND_net), 
            .\dc32_fifo_data_out[5] (dc32_fifo_data_out[5]), .\dc32_fifo_data_out[4] (dc32_fifo_data_out[4]), 
            .\dc32_fifo_data_out[3] (dc32_fifo_data_out[3]), .\dc32_fifo_data_out[2] (dc32_fifo_data_out[2]), 
            .\dc32_fifo_data_out[1] (dc32_fifo_data_out[1]), .DEBUG_5_c_0(DEBUG_5_c_0), 
            .DEBUG_2_c(DEBUG_2_c), .sc32_fifo_read_enable(sc32_fifo_read_enable), 
            .n5367(n5367), .n5366(n5366), .n5365(n5365), .n5364(n5364), 
            .n5363(n5363), .n5362(n5362), .n5361(n5361), .n5360(n5360), 
            .n5359(n5359), .n5358(n5358), .n5357(n5357), .n5356(n5356), 
            .n5355(n5355), .n5354(n5354), .n5353(n5353), .n5352(n5352), 
            .n5351(n5351), .n5350(n5350), .n5349(n5349), .n5348(n5348), 
            .n5347(n5347), .n5346(n5346), .n5345(n5345), .n5344(n5344), 
            .n5343(n5343), .n5342(n5342), .n5341(n5341), .n5340(n5340), 
            .n5339(n5339), .n5338(n5338), .n5337(n5337)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(620[20] 634[2])
    SB_LUT4 i5494_2_lut_3_lut (.I0(DEBUG_9_c_0), .I1(bluejay_data_out_31__N_921), 
            .I2(bluejay_data_out_31__N_922), .I3(GND_net), .O(n6968));   // src/bluejay_data.v(134[8] 156[4])
    defparam i5494_2_lut_3_lut.LUT_INIT = 16'ha8a8;
    \uart_tx(CLKS_PER_BIT=20)  pc_tx (.GND_net(GND_net), .VCC_net(VCC_net), 
            .UART_TX_c(UART_TX_c), .SLM_CLK_c(SLM_CLK_c), .r_SM_Main({r_SM_Main_adj_1467}), 
            .\r_SM_Main_2__N_1026[1] (r_SM_Main_2__N_1026[1]), .\r_Bit_Index[0] (r_Bit_Index_adj_1469[0]), 
            .n6966(n6966), .r_Tx_Data({r_Tx_Data}), .n6965(n6965), .n6964(n6964), 
            .n6963(n6963), .n6962(n6962), .n6961(n6961), .n6960(n6960), 
            .n6950(n6950), .n16231(n16231), .n5024(n5024), .n5460(n5460), 
            .\r_SM_Main_2__N_1029[0] (r_SM_Main_2__N_1029[0]), .n4314(n4314), 
            .n5576(n5576), .n5575(n5575), .tx_uart_active_flag(tx_uart_active_flag), 
            .n4(n4_adj_1442)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(859[42] 868[3])
    SB_LUT4 i3910_1_lut_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n5384));   // src/top.v(1165[8] 1232[4])
    defparam i3910_1_lut_2_lut.LUT_INIT = 16'h7777;
    usb3_if usb3_if_inst (.reset_per_frame(reset_per_frame), .reset_per_frame_latched(reset_per_frame_latched), 
            .SLM_CLK_c(SLM_CLK_c), .dc32_fifo_empty(dc32_fifo_empty), .VCC_net(VCC_net), 
            .FT_RD_c(FT_RD_c), .FIFO_CLK_c(FIFO_CLK_c), .dc32_fifo_data_in({dc32_fifo_data_in}), 
            .dc32_fifo_write_enable(dc32_fifo_write_enable), .buffer_switch_done(buffer_switch_done), 
            .buffer_switch_done_latched(buffer_switch_done_latched), .GND_net(GND_net), 
            .DEBUG_1_c(DEBUG_1_c), .n663(n663), .n7014(n7014), .FR_RXF_c(FR_RXF_c), 
            .FT_OE_c(FT_OE_c), .DEBUG_3_c_0_c(DEBUG_3_c_0_c), .FIFO_D1_c_1(FIFO_D1_c_1), 
            .FIFO_D2_c_2(FIFO_D2_c_2), .FIFO_D3_c_3(FIFO_D3_c_3), .FIFO_D4_c_4(FIFO_D4_c_4), 
            .FIFO_D5_c_5(FIFO_D5_c_5), .FIFO_D6_c_6(FIFO_D6_c_6), .FIFO_D7_c_7(FIFO_D7_c_7), 
            .FIFO_D8_c_8(FIFO_D8_c_8), .FIFO_D9_c_9(FIFO_D9_c_9), .FIFO_D10_c_10(FIFO_D10_c_10), 
            .FIFO_D11_c_11(FIFO_D11_c_11), .FIFO_D12_c_12(FIFO_D12_c_12), 
            .FIFO_D13_c_13(FIFO_D13_c_13), .FIFO_D14_c_14(FIFO_D14_c_14), 
            .FIFO_D15_c_15(FIFO_D15_c_15), .FIFO_D16_c_16(FIFO_D16_c_16), 
            .FIFO_D17_c_17(FIFO_D17_c_17), .FIFO_D18_c_18(FIFO_D18_c_18), 
            .FIFO_D19_c_19(FIFO_D19_c_19), .FIFO_D20_c_20(FIFO_D20_c_20), 
            .FIFO_D21_c_21(FIFO_D21_c_21), .FIFO_D22_c_22(FIFO_D22_c_22), 
            .FIFO_D23_c_23(FIFO_D23_c_23), .FIFO_D24_c_24(FIFO_D24_c_24), 
            .FIFO_D25_c_25(FIFO_D25_c_25), .FIFO_D26_c_26(FIFO_D26_c_26), 
            .FIFO_D27_c_27(FIFO_D27_c_27), .FIFO_D28_c_28(FIFO_D28_c_28), 
            .FIFO_D29_c_29(FIFO_D29_c_29), .FIFO_D30_c_30(FIFO_D30_c_30), 
            .FIFO_D31_c_31(FIFO_D31_c_31)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(544[9] 560[3])
    clock clock_inst (.GND_net(GND_net), .VCC_net(VCC_net), .ICE_SYSCLK_c(ICE_SYSCLK_c), 
          .pll_clk_unbuf(pll_clk_unbuf)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(222[7] 228[3])
    spi spi0 (.n4837(n4837), .SLM_CLK_c(SLM_CLK_c), .GND_net(GND_net), 
        .tx_addr_byte({tx_addr_byte}), .n2407(n2407), .SEN_c_1(SEN_c_1), 
        .\tx_data_byte[7] (tx_data_byte[7]), .SOUT_c(SOUT_c), .n4884(n4884), 
        .\rx_shift_reg[0] (rx_shift_reg[0]), .SDAT_c_15(SDAT_c_15), .n6988(n6988), 
        .rx_buf_byte({rx_buf_byte}), .n6987(n6987), .n6986(n6986), .n6985(n6985), 
        .n6984(n6984), .n6983(n6983), .n6982(n6982), .n6981(n6981), 
        .\rx_shift_reg[7] (rx_shift_reg[7]), .n6980(n6980), .\rx_shift_reg[6] (rx_shift_reg[6]), 
        .n6979(n6979), .\rx_shift_reg[5] (rx_shift_reg[5]), .n6978(n6978), 
        .\rx_shift_reg[4] (rx_shift_reg[4]), .n6977(n6977), .\rx_shift_reg[3] (rx_shift_reg[3]), 
        .n6976(n6976), .\rx_shift_reg[2] (rx_shift_reg[2]), .n6975(n6975), 
        .\rx_shift_reg[1] (rx_shift_reg[1]), .n12537(n12537), .VCC_net(VCC_net), 
        .\tx_shift_reg[0] (tx_shift_reg[0]), .\tx_data_byte[1] (tx_data_byte[1]), 
        .multi_byte_spi_trans_flag_r(multi_byte_spi_trans_flag_r), .\tx_data_byte[2] (tx_data_byte[2]), 
        .\tx_data_byte[3] (tx_data_byte[3]), .\tx_data_byte[4] (tx_data_byte[4]), 
        .spi_rx_byte_ready(spi_rx_byte_ready), .SCK_c_0(SCK_c_0), .spi_start_transfer_r(spi_start_transfer_r), 
        .n5578(n5578), .\tx_data_byte[5] (tx_data_byte[5]), .\tx_data_byte[6] (tx_data_byte[6]), 
        .n3963(n3963)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(924[5] 948[2])
>>>>>>> master
    
endmodule
//
// Verilog Description of module timing_controller
//

<<<<<<< HEAD
module timing_controller (SLM_CLK_c, GND_net, sc32_fifo_read_enable, n10668, 
            VCC_net, state, dc32_fifo_read_enable, n1967, DEBUG_8_c, 
            DEBUG_6_c, n63, n5132, \state_timeout_counter[7] , n3, 
            n11094, n5500, n1459, n106, n80, n5504, buffer_switch_done, 
            n2072, n7836, INVERT_c_4, n11257, dc32_fifo_full, n11101, 
            n7, n59, n6, \aempty_flag_impl.ae_flag_nxt_w , n4943, 
            n47, reset_all, n11700, reset_per_frame, n8057, line_of_data_available, 
            UPDATE_c_3) /* synthesis syn_module_defined=1 */ ;
    input SLM_CLK_c;
    input GND_net;
    output sc32_fifo_read_enable;
    input n10668;
    input VCC_net;
    output [3:0]state;
    output dc32_fifo_read_enable;
    input n1967;
    input DEBUG_8_c;
    input DEBUG_6_c;
    output n63;
    output n5132;
    input \state_timeout_counter[7] ;
    input n3;
    input n11094;
    output n5500;
    input n1459;
    input n106;
    input n80;
    output n5504;
    output buffer_switch_done;
    input n2072;
    input n7836;
    output INVERT_c_4;
    output n11257;
    input dc32_fifo_full;
    output n11101;
    input n7;
    input n59;
    input n6;
    output \aempty_flag_impl.ae_flag_nxt_w ;
    output n4943;
    output n47;
    output reset_all;
    input n11700;
    output reset_per_frame;
    input n8057;
    output line_of_data_available;
    output UPDATE_c_3;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [31:0]n2145;
    
    wire n5068;
    wire [31:0]state_timeout_counter;   // src/timing_controller.v(80[12:33])
    wire [31:0]n630;
    
    wire n5537, n11156, n6461;
    wire [2:0]fifo_state;   // src/timing_controller.v(77[11:21])
    
    wire n40, sc32_fifo_read_enable_N_366;
    wire [2:0]fifo_state_2__N_80;
    
    wire n23;
    wire [3:0]state_3__N_83;
    
    wire n11119, dc32_fifo_read_enable_N_359, n11406, n10274, n10275, 
        n10253, n10254, n11382, n10252, n7264, n11049, n11050, 
        n4070, n6520, n3_c, n69, n4, n31, n7261, n10273, n7265, 
        n7269, n8067, n10393;
    wire [5:0]fifo_state_timeout_counter;   // src/timing_controller.v(79[11:37])
    
    wire n10295, n4_adj_1391, n7_c, n10272;
    wire [6:0]fifo_state_timeout_counter_5__N_125;
    
    wire n10294, n10293, n5, n10292, n11118, n10271, n10291, n11352, 
        n26, n10676, n11379;
    wire [31:0]n2073;
    
    wire n2106, n2144, n11347, n11378, n11092, n11377, n11376, 
        n11375, n11374, n11373, n4068, n10270, n11191, n10251, 
        n10269, n10268, n10267, n10266, n10250;
    wire [4:0]n1103;
    
    wire n4_adj_1392, n11358, n10265, n5304, n10264, n10263, n10262, 
        n11356, n10261, n10260, n10259, n38, n52, n5496, n56, 
        n54, n55, n11102, n28, n10258, n10, n53, n50, n10257, 
        n58, n62, n49, n10280, n10279, n10278, n11506, n2, n10277, 
        n10256, n10276, n11104, n10255, n11391;
    
    SB_DFFE state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(SLM_CLK_c), 
            .E(n5068), .D(n2145[0]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i22 (.Q(state_timeout_counter[22]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[22]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 i41_3_lut (.I0(n11156), .I1(n6461), .I2(fifo_state[0]), .I3(GND_net), 
            .O(n40));   // src/timing_controller.v(78[11:16])
    defparam i41_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF sc32_fifo_read_enable_92 (.Q(sc32_fifo_read_enable), .C(SLM_CLK_c), 
           .D(sc32_fifo_read_enable_N_366));   // src/timing_controller.v(88[8] 151[4])
    SB_DFFE fifo_state_i0 (.Q(fifo_state[0]), .C(SLM_CLK_c), .E(n23), 
            .D(fifo_state_2__N_80[0]));   // src/timing_controller.v(88[8] 151[4])
    SB_DFFE state_i3 (.Q(state[3]), .C(SLM_CLK_c), .E(VCC_net), .D(n10668));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_i0 (.Q(state[0]), .C(SLM_CLK_c), .E(n11119), .D(state_3__N_83[0]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFF dc32_fifo_read_enable_90 (.Q(dc32_fifo_read_enable), .C(SLM_CLK_c), 
           .D(dc32_fifo_read_enable_N_359));   // src/timing_controller.v(88[8] 151[4])
    SB_LUT4 i9912_2_lut (.I0(fifo_state[0]), .I1(n6461), .I2(GND_net), 
            .I3(GND_net), .O(n11406));   // src/timing_controller.v(93[5] 150[12])
    defparam i9912_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY sub_71_add_2_27 (.CI(n10274), .I0(state_timeout_counter[25]), 
            .I1(VCC_net), .CO(n10275));
    SB_CARRY sub_71_add_2_6 (.CI(n10253), .I0(state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n10254));
    SB_LUT4 sub_71_add_2_5_lut (.I0(n1967), .I1(state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n10252), .O(n11382)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_5_lut.LUT_INIT = 16'h8228;
=======
module timing_controller (SLM_CLK_c, DEBUG_2_c, sc32_fifo_read_enable, 
            state, dc32_fifo_read_enable, n63, GND_net, VCC_net, n2075, 
            n2180, n9015, buffer_switch_done, n12477, n8659, reset_all, 
            line_of_data_available, n7, n8, \aempty_flag_impl.ae_flag_nxt_w , 
            INVERT_c_4, n4903, get_next_word, dc32_fifo_almost_empty, 
            n4688, dc32_fifo_full, n9013, n12884, reset_per_frame, 
            UPDATE_c_3, n25, n12882) /* synthesis syn_module_defined=1 */ ;
    input SLM_CLK_c;
    output DEBUG_2_c;
    output sc32_fifo_read_enable;
    output [3:0]state;
    output dc32_fifo_read_enable;
    output n63;
    input GND_net;
    input VCC_net;
    input n2075;
    input n2180;
    output n9015;
    output buffer_switch_done;
    input n12477;
    input n8659;
    output reset_all;
    output line_of_data_available;
    input n7;
    input n8;
    output \aempty_flag_impl.ae_flag_nxt_w ;
    output INVERT_c_4;
    output n4903;
    input get_next_word;
    input dc32_fifo_almost_empty;
    input n4688;
    input dc32_fifo_full;
    input n9013;
    input n12884;
    output reset_per_frame;
    output UPDATE_c_3;
    output n25;
    output n12882;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n12866, n8325;
    wire [5:0]fifo_state_timeout_counter;   // src/timing_controller.v(79[11:37])
    
    wire n11540;
    wire [31:0]n2253;
    
    wire n4838;
    wire [31:0]state_timeout_counter;   // src/timing_controller.v(80[12:33])
    
    wire sc32_fifo_write_enable_N_366, sc32_fifo_read_enable_N_367;
    wire [2:0]fifo_state_2__N_80;
    
    wire n13044;
    wire [2:0]fifo_state;   // src/timing_controller.v(77[11:21])
    wire [6:0]fifo_state_timeout_counter_5__N_125;
    
    wire n8321, n12868;
    wire [3:0]state_3__N_83;
    
    wire n12908, dc32_fifo_read_enable_N_359, n2334, n14260, n12074, 
        n12089, n12090, n14282;
    wire [31:0]n2181;
    
    wire n2252, n14279, n9023, n14283, n14284, n14285, n14286, 
        n12902, n14287, n14288, n14289, n14290, n14291, n14292, 
        n14293, n1290, n11566, n14255, n18, n12499, n4, n14281, 
        n14280, n12893;
    wire [4:0]n1138;
    
    wire n12075, n12088, n12073, n12072;
    wire [31:0]n628;
    
    wire n12087, n5419, n5404, n12086, n12914, n12085, n4936, 
        n12084, n12071, n12083, n14248, n12101, n12100, n12099, 
        n12082, n12098, n12865, n12126, n94, n12081, n12125, n12097, 
        n12096, n12095, n12080, n12124, n12079, n12078, n12123, 
        n12094, n12093, n12122, n12092, n12077, n12883, n12076, 
        n2, n8043, n14311, n16, n7_adj_1412, n7_adj_1413, n15, 
        n12988, n70, n96, n14276, n11, n12091, n5, n38, n52, 
        n56, n54, n55, n53, n50, n58, n62, n49, n14398, n17, 
        n12900, n4_adj_1414;
    
    SB_DFFESS fifo_state_timeout_counter_i0_i5 (.Q(fifo_state_timeout_counter[5]), 
            .C(SLM_CLK_c), .E(n8325), .D(n12866), .S(n11540));   // src/timing_controller.v(88[8] 151[4])
    SB_DFFE state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2253[0]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFF sc32_fifo_write_enable_89 (.Q(DEBUG_2_c), .C(SLM_CLK_c), .D(sc32_fifo_write_enable_N_366));   // src/timing_controller.v(88[8] 151[4])
    SB_DFF sc32_fifo_read_enable_90 (.Q(sc32_fifo_read_enable), .C(SLM_CLK_c), 
           .D(sc32_fifo_read_enable_N_367));   // src/timing_controller.v(88[8] 151[4])
    SB_DFFE fifo_state_i0 (.Q(fifo_state[0]), .C(SLM_CLK_c), .E(n13044), 
            .D(fifo_state_2__N_80[0]));   // src/timing_controller.v(88[8] 151[4])
    SB_DFFESR fifo_state_timeout_counter_i0_i4 (.Q(fifo_state_timeout_counter[4]), 
            .C(SLM_CLK_c), .E(n8325), .D(fifo_state_timeout_counter_5__N_125[4]), 
            .R(n8321));   // src/timing_controller.v(88[8] 151[4])
    SB_DFFESR fifo_state_timeout_counter_i0_i3 (.Q(fifo_state_timeout_counter[3]), 
            .C(SLM_CLK_c), .E(n8325), .D(n12868), .R(n11540));   // src/timing_controller.v(88[8] 151[4])
    SB_DFFE state_i0 (.Q(state[0]), .C(SLM_CLK_c), .E(n12908), .D(state_3__N_83[0]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFF dc32_fifo_read_enable_88 (.Q(dc32_fifo_read_enable), .C(SLM_CLK_c), 
           .D(dc32_fifo_read_enable_N_359));   // src/timing_controller.v(88[8] 151[4])
    SB_DFFESR fifo_state_timeout_counter_i0_i2 (.Q(fifo_state_timeout_counter[2]), 
            .C(SLM_CLK_c), .E(n8325), .D(fifo_state_timeout_counter_5__N_125[2]), 
            .R(n8321));   // src/timing_controller.v(88[8] 151[4])
    SB_DFFESR fifo_state_timeout_counter_i0_i1 (.Q(fifo_state_timeout_counter[1]), 
            .C(SLM_CLK_c), .E(n8325), .D(fifo_state_timeout_counter_5__N_125[1]), 
            .R(n8321));   // src/timing_controller.v(88[8] 151[4])
    SB_LUT4 state_3__I_0_103_Mux_2_i15_4_lut (.I0(state[1]), .I1(state[2]), 
            .I2(state[3]), .I3(state[0]), .O(state_3__N_83[2]));   // src/timing_controller.v(160[5] 229[12])
    defparam state_3__I_0_103_Mux_2_i15_4_lut.LUT_INIT = 16'hc2ce;
    SB_LUT4 i1113_2_lut_3_lut (.I0(state[0]), .I1(n63), .I2(state[1]), 
            .I3(GND_net), .O(n2334));   // src/timing_controller.v(154[8] 230[4])
    defparam i1113_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 sub_69_add_2_6_lut (.I0(n2075), .I1(state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n12074), .O(n14260)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_69_add_2_21 (.CI(n12089), .I0(state_timeout_counter[19]), 
            .I1(VCC_net), .CO(n12090));
    SB_LUT4 mux_1055_i4_3_lut (.I0(n14282), .I1(state[1]), .I2(n2180), 
            .I3(GND_net), .O(n2181[3]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1055_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10875_4_lut (.I0(n14260), .I1(state[1]), .I2(n2180), .I3(n2252), 
            .O(n2253[4]));   // src/timing_controller.v(160[5] 229[12])
    defparam i10875_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_1063_i6_3_lut (.I0(n14279), .I1(state[1]), .I2(n2252), 
            .I3(GND_net), .O(n2253[5]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1063_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7554_2_lut_3_lut (.I0(state[1]), .I1(state[2]), .I2(n63), 
            .I3(GND_net), .O(n9023));
    defparam i7554_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i7546_2_lut_3_lut (.I0(state[1]), .I1(state[2]), .I2(state[0]), 
            .I3(GND_net), .O(n9015));
    defparam i7546_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_1055_i10_3_lut (.I0(n14283), .I1(state[1]), .I2(n2180), 
            .I3(GND_net), .O(n2181[9]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1055_i10_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1055_i11_3_lut (.I0(n14284), .I1(state[1]), .I2(n2180), 
            .I3(GND_net), .O(n2181[10]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1055_i11_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1055_i13_3_lut (.I0(n14285), .I1(state[1]), .I2(n2180), 
            .I3(GND_net), .O(n2181[12]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1055_i13_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1055_i15_3_lut (.I0(n14286), .I1(state[1]), .I2(n2180), 
            .I3(GND_net), .O(n2181[14]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1055_i15_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1063_i4_3_lut_4_lut (.I0(state[1]), .I1(n12902), .I2(n2252), 
            .I3(n2181[3]), .O(n2253[3]));   // src/timing_controller.v(154[8] 230[4])
    defparam mux_1063_i4_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_1055_i16_3_lut (.I0(n14287), .I1(state[1]), .I2(n2180), 
            .I3(GND_net), .O(n2181[15]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1055_i16_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1055_i19_3_lut (.I0(n14288), .I1(state[1]), .I2(n2180), 
            .I3(GND_net), .O(n2181[18]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1055_i19_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1055_i20_3_lut (.I0(n14289), .I1(state[1]), .I2(n2180), 
            .I3(GND_net), .O(n2181[19]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1055_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1063_i10_3_lut_4_lut (.I0(state[1]), .I1(n12902), .I2(n2252), 
            .I3(n2181[9]), .O(n2253[9]));   // src/timing_controller.v(154[8] 230[4])
    defparam mux_1063_i10_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_1063_i11_3_lut_4_lut (.I0(state[1]), .I1(n12902), .I2(n2252), 
            .I3(n2181[10]), .O(n2253[10]));   // src/timing_controller.v(154[8] 230[4])
    defparam mux_1063_i11_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_1055_i21_3_lut (.I0(n14290), .I1(state[1]), .I2(n2180), 
            .I3(GND_net), .O(n2181[20]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1055_i21_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1055_i23_3_lut (.I0(n14291), .I1(state[1]), .I2(n2180), 
            .I3(GND_net), .O(n2181[22]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1055_i23_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1055_i24_3_lut (.I0(n14292), .I1(state[1]), .I2(n2180), 
            .I3(GND_net), .O(n2181[23]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1055_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1063_i13_3_lut_4_lut (.I0(state[1]), .I1(n12902), .I2(n2252), 
            .I3(n2181[12]), .O(n2253[12]));   // src/timing_controller.v(154[8] 230[4])
    defparam mux_1063_i13_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_1055_i25_3_lut (.I0(n14293), .I1(state[1]), .I2(n2180), 
            .I3(GND_net), .O(n2181[24]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1055_i25_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1063_i15_3_lut_4_lut (.I0(state[1]), .I1(n12902), .I2(n2252), 
            .I3(n2181[14]), .O(n2253[14]));   // src/timing_controller.v(154[8] 230[4])
    defparam mux_1063_i15_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_1063_i16_3_lut_4_lut (.I0(state[1]), .I1(n12902), .I2(n2252), 
            .I3(n2181[15]), .O(n2253[15]));   // src/timing_controller.v(154[8] 230[4])
    defparam mux_1063_i16_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_1063_i19_3_lut_4_lut (.I0(state[1]), .I1(n12902), .I2(n2252), 
            .I3(n2181[18]), .O(n2253[18]));   // src/timing_controller.v(154[8] 230[4])
    defparam mux_1063_i19_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 i12265_3_lut (.I0(fifo_state[1]), .I1(fifo_state[0]), .I2(fifo_state[2]), 
            .I3(GND_net), .O(fifo_state_2__N_80[1]));   // src/timing_controller.v(93[5] 150[12])
    defparam i12265_3_lut.LUT_INIT = 16'ha6a6;
    SB_LUT4 i12220_4_lut (.I0(n1290), .I1(n11566), .I2(fifo_state[0]), 
            .I3(fifo_state[2]), .O(n14255));
    defparam i12220_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36_4_lut (.I0(n14255), .I1(n18), .I2(fifo_state[1]), .I3(fifo_state[2]), 
            .O(n12499));
    defparam i36_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_1063_i20_3_lut_4_lut (.I0(state[1]), .I1(n12902), .I2(n2252), 
            .I3(n2181[19]), .O(n2253[19]));   // src/timing_controller.v(154[8] 230[4])
    defparam mux_1063_i20_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_1063_i21_3_lut_4_lut (.I0(state[1]), .I1(n12902), .I2(n2252), 
            .I3(n2181[20]), .O(n2253[20]));   // src/timing_controller.v(154[8] 230[4])
    defparam mux_1063_i21_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 i12_3_lut (.I0(fifo_state[1]), .I1(fifo_state[2]), .I2(fifo_state[0]), 
            .I3(GND_net), .O(fifo_state_2__N_80[2]));   // src/timing_controller.v(77[11:21])
    defparam i12_3_lut.LUT_INIT = 16'h2c2c;
    SB_LUT4 i1_2_lut (.I0(n2075), .I1(n2180), .I2(GND_net), .I3(GND_net), 
            .O(n4));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_1055_i3_3_lut (.I0(n14281), .I1(state[1]), .I2(n2180), 
            .I3(GND_net), .O(n2181[2]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1055_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1055_i2_3_lut (.I0(n14280), .I1(state[1]), .I2(n2180), 
            .I3(GND_net), .O(n2181[1]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1055_i2_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1063_i25_3_lut_4_lut (.I0(state[1]), .I1(n12902), .I2(n2252), 
            .I3(n2181[24]), .O(n2253[24]));   // src/timing_controller.v(154[8] 230[4])
    defparam mux_1063_i25_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(state[1]), .I1(state[3]), .I2(state[2]), 
            .I3(state[0]), .O(n12893));   // src/timing_controller.v(160[5] 229[12])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 mux_1063_i24_3_lut_4_lut (.I0(state[1]), .I1(n12902), .I2(n2252), 
            .I3(n2181[23]), .O(n2253[23]));   // src/timing_controller.v(154[8] 230[4])
    defparam mux_1063_i24_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_1063_i23_3_lut_4_lut (.I0(state[1]), .I1(n12902), .I2(n2252), 
            .I3(n2181[22]), .O(n2253[22]));   // src/timing_controller.v(154[8] 230[4])
    defparam mux_1063_i23_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_DFF invert_98_i2 (.Q(buffer_switch_done), .C(SLM_CLK_c), .D(n12893));   // src/timing_controller.v(160[5] 229[12])
    SB_DFFE state_i3 (.Q(state[3]), .C(SLM_CLK_c), .E(VCC_net), .D(n12477));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 mux_379_Mux_4_i15_4_lut_4_lut (.I0(state[2]), .I1(state[0]), 
            .I2(state[1]), .I3(state[3]), .O(n1138[4]));
    defparam mux_379_Mux_4_i15_4_lut_4_lut.LUT_INIT = 16'h01a0;
    SB_CARRY sub_69_add_2_6 (.CI(n12074), .I0(state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n12075));
    SB_LUT4 sub_69_add_2_20_lut (.I0(n2075), .I1(state_timeout_counter[18]), 
            .I2(VCC_net), .I3(n12088), .O(n14288)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_69_add_2_5_lut (.I0(n2075), .I1(state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n12073), .O(n14282)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_69_add_2_5 (.CI(n12073), .I0(state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n12074));
    SB_CARRY sub_69_add_2_20 (.CI(n12088), .I0(state_timeout_counter[18]), 
            .I1(VCC_net), .CO(n12089));
    SB_LUT4 sub_69_add_2_4_lut (.I0(n8659), .I1(state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n12072), .O(n14281)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_69_add_2_19_lut (.I0(GND_net), .I1(state_timeout_counter[17]), 
            .I2(VCC_net), .I3(n12087), .O(n628[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_19 (.CI(n12087), .I0(state_timeout_counter[17]), 
            .I1(VCC_net), .CO(n12088));
    SB_DFFESR state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2181[1]), .R(n5419));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2181[2]), .R(n5419));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i6 (.Q(state_timeout_counter[6]), .C(SLM_CLK_c), 
            .E(n4838), .D(n628[6]), .R(n5404));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i7 (.Q(state_timeout_counter[7]), .C(SLM_CLK_c), 
            .E(n4838), .D(n628[7]), .R(n5404));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i8 (.Q(state_timeout_counter[8]), .C(SLM_CLK_c), 
            .E(n4838), .D(n628[8]), .R(n5404));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE fifo_state_i2 (.Q(fifo_state[2]), .C(SLM_CLK_c), .E(n12499), 
            .D(fifo_state_2__N_80[2]));   // src/timing_controller.v(88[8] 151[4])
    SB_DFFESR state_timeout_counter_i0_i11 (.Q(state_timeout_counter[11]), 
            .C(SLM_CLK_c), .E(n4838), .D(n628[11]), .R(n5404));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i13 (.Q(state_timeout_counter[13]), 
            .C(SLM_CLK_c), .E(n4838), .D(n628[13]), .R(n5404));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i16 (.Q(state_timeout_counter[16]), 
            .C(SLM_CLK_c), .E(n4838), .D(n628[16]), .R(n5404));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i17 (.Q(state_timeout_counter[17]), 
            .C(SLM_CLK_c), .E(n4838), .D(n628[17]), .R(n5404));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 sub_69_add_2_18_lut (.I0(GND_net), .I1(state_timeout_counter[16]), 
            .I2(VCC_net), .I3(n12086), .O(n628[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR state_timeout_counter_i0_i21 (.Q(state_timeout_counter[21]), 
            .C(SLM_CLK_c), .E(n4838), .D(n628[21]), .R(n5404));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i25 (.Q(state_timeout_counter[25]), 
            .C(SLM_CLK_c), .E(n4838), .D(n628[25]), .R(n5404));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i26 (.Q(state_timeout_counter[26]), 
            .C(SLM_CLK_c), .E(n4838), .D(n628[26]), .R(n5404));   // src/timing_controller.v(154[8] 230[4])
    SB_CARRY sub_69_add_2_4 (.CI(n12072), .I0(state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n12073));
    SB_DFFESR state_timeout_counter_i0_i27 (.Q(state_timeout_counter[27]), 
            .C(SLM_CLK_c), .E(n4838), .D(n628[27]), .R(n5404));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i28 (.Q(state_timeout_counter[28]), 
            .C(SLM_CLK_c), .E(n4838), .D(n628[28]), .R(n5404));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i29 (.Q(state_timeout_counter[29]), 
            .C(SLM_CLK_c), .E(n4838), .D(n628[29]), .R(n5404));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i30 (.Q(state_timeout_counter[30]), 
            .C(SLM_CLK_c), .E(n4838), .D(n628[30]), .R(n5404));   // src/timing_controller.v(154[8] 230[4])
    SB_CARRY sub_69_add_2_18 (.CI(n12086), .I0(state_timeout_counter[16]), 
            .I1(VCC_net), .CO(n12087));
    SB_DFFESR state_timeout_counter_i0_i31 (.Q(state_timeout_counter[31]), 
            .C(SLM_CLK_c), .E(n4838), .D(n628[31]), .R(n5404));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE fifo_state_i1 (.Q(fifo_state[1]), .C(SLM_CLK_c), .E(n13044), 
            .D(fifo_state_2__N_80[1]));   // src/timing_controller.v(88[8] 151[4])
    SB_LUT4 i1_2_lut_3_lut (.I0(state[2]), .I1(state[0]), .I2(n63), .I3(GND_net), 
            .O(n12914));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_DFFE state_timeout_counter_i0_i24 (.Q(state_timeout_counter[24]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2253[24]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i23 (.Q(state_timeout_counter[23]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2253[23]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i22 (.Q(state_timeout_counter[22]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2253[22]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i20 (.Q(state_timeout_counter[20]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2253[20]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i19 (.Q(state_timeout_counter[19]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2253[19]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i18 (.Q(state_timeout_counter[18]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2253[18]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i15 (.Q(state_timeout_counter[15]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2253[15]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i14 (.Q(state_timeout_counter[14]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2253[14]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i12 (.Q(state_timeout_counter[12]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2253[12]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i10 (.Q(state_timeout_counter[10]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2253[10]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i9 (.Q(state_timeout_counter[9]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2253[9]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i5 (.Q(state_timeout_counter[5]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2253[5]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2253[4]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(SLM_CLK_c), 
            .E(n4838), .D(n2253[3]));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 sub_69_add_2_17_lut (.I0(n2075), .I1(state_timeout_counter[15]), 
            .I2(VCC_net), .I3(n12085), .O(n14287)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_69_add_2_17 (.CI(n12085), .I0(state_timeout_counter[15]), 
            .I1(VCC_net), .CO(n12086));
    SB_DFFE state_i1 (.Q(state[1]), .C(SLM_CLK_c), .E(n4936), .D(state_3__N_83[1]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_i2 (.Q(state[2]), .C(SLM_CLK_c), .E(n4936), .D(state_3__N_83[2]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR fifo_state_timeout_counter_i0_i0 (.Q(fifo_state_timeout_counter[0]), 
            .C(SLM_CLK_c), .E(n8325), .D(fifo_state_timeout_counter_5__N_125[0]), 
            .R(n8321));   // src/timing_controller.v(88[8] 151[4])
    SB_LUT4 sub_69_add_2_16_lut (.I0(n2075), .I1(state_timeout_counter[14]), 
            .I2(VCC_net), .I3(n12084), .O(n14286)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_69_add_2_3_lut (.I0(n2075), .I1(state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n12071), .O(n14280)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_69_add_2_16 (.CI(n12084), .I0(state_timeout_counter[14]), 
            .I1(VCC_net), .CO(n12085));
    SB_LUT4 sub_69_add_2_15_lut (.I0(GND_net), .I1(state_timeout_counter[13]), 
            .I2(VCC_net), .I3(n12083), .O(n628[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_3 (.CI(n12071), .I0(state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n12072));
    SB_LUT4 sub_69_add_2_2_lut (.I0(n8659), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n14248)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_69_add_2_2 (.CI(VCC_net), .I0(state_timeout_counter[0]), 
            .I1(GND_net), .CO(n12071));
    SB_LUT4 sub_69_add_2_33_lut (.I0(GND_net), .I1(state_timeout_counter[31]), 
            .I2(VCC_net), .I3(n12101), .O(n628[31])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_69_add_2_32_lut (.I0(GND_net), .I1(state_timeout_counter[30]), 
            .I2(VCC_net), .I3(n12100), .O(n628[30])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_32 (.CI(n12100), .I0(state_timeout_counter[30]), 
            .I1(VCC_net), .CO(n12101));
    SB_CARRY sub_69_add_2_15 (.CI(n12083), .I0(state_timeout_counter[13]), 
            .I1(VCC_net), .CO(n12084));
    SB_LUT4 sub_69_add_2_31_lut (.I0(GND_net), .I1(state_timeout_counter[29]), 
            .I2(VCC_net), .I3(n12099), .O(n628[29])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_69_add_2_14_lut (.I0(n2075), .I1(state_timeout_counter[12]), 
            .I2(VCC_net), .I3(n12082), .O(n14285)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_69_add_2_31 (.CI(n12099), .I0(state_timeout_counter[29]), 
            .I1(VCC_net), .CO(n12100));
    SB_LUT4 sub_69_add_2_30_lut (.I0(GND_net), .I1(state_timeout_counter[28]), 
            .I2(VCC_net), .I3(n12098), .O(n628[28])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_14 (.CI(n12082), .I0(state_timeout_counter[12]), 
            .I1(VCC_net), .CO(n12083));
    SB_LUT4 sub_111_add_2_7_lut (.I0(n94), .I1(fifo_state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n12126), .O(n12865)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_69_add_2_13_lut (.I0(GND_net), .I1(state_timeout_counter[11]), 
            .I2(VCC_net), .I3(n12081), .O(n628[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_30 (.CI(n12098), .I0(state_timeout_counter[28]), 
            .I1(VCC_net), .CO(n12099));
    SB_LUT4 sub_111_add_2_6_lut (.I0(GND_net), .I1(fifo_state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n12125), .O(fifo_state_timeout_counter_5__N_125[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_69_add_2_29_lut (.I0(GND_net), .I1(state_timeout_counter[27]), 
            .I2(VCC_net), .I3(n12097), .O(n628[27])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_111_add_2_6 (.CI(n12125), .I0(fifo_state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n12126));
    SB_CARRY sub_69_add_2_29 (.CI(n12097), .I0(state_timeout_counter[27]), 
            .I1(VCC_net), .CO(n12098));
    SB_LUT4 sub_69_add_2_28_lut (.I0(GND_net), .I1(state_timeout_counter[26]), 
            .I2(VCC_net), .I3(n12096), .O(n628[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_13 (.CI(n12081), .I0(state_timeout_counter[11]), 
            .I1(VCC_net), .CO(n12082));
    SB_CARRY sub_69_add_2_28 (.CI(n12096), .I0(state_timeout_counter[26]), 
            .I1(VCC_net), .CO(n12097));
    SB_LUT4 sub_69_add_2_27_lut (.I0(GND_net), .I1(state_timeout_counter[25]), 
            .I2(VCC_net), .I3(n12095), .O(n628[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_69_add_2_12_lut (.I0(n2075), .I1(state_timeout_counter[10]), 
            .I2(VCC_net), .I3(n12080), .O(n14284)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_111_add_2_5_lut (.I0(GND_net), .I1(fifo_state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n12124), .O(fifo_state_timeout_counter_5__N_125[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_12 (.CI(n12080), .I0(state_timeout_counter[10]), 
            .I1(VCC_net), .CO(n12081));
    SB_LUT4 sub_69_add_2_11_lut (.I0(n2075), .I1(state_timeout_counter[9]), 
            .I2(VCC_net), .I3(n12079), .O(n14283)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_111_add_2_5 (.CI(n12124), .I0(fifo_state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n12125));
    SB_CARRY sub_69_add_2_11 (.CI(n12079), .I0(state_timeout_counter[9]), 
            .I1(VCC_net), .CO(n12080));
    SB_CARRY sub_69_add_2_27 (.CI(n12095), .I0(state_timeout_counter[25]), 
            .I1(VCC_net), .CO(n12096));
    SB_LUT4 sub_69_add_2_10_lut (.I0(GND_net), .I1(state_timeout_counter[8]), 
            .I2(VCC_net), .I3(n12078), .O(n628[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_111_add_2_4_lut (.I0(GND_net), .I1(fifo_state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n12123), .O(fifo_state_timeout_counter_5__N_125[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_69_add_2_26_lut (.I0(n2075), .I1(state_timeout_counter[24]), 
            .I2(VCC_net), .I3(n12094), .O(n14293)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_69_add_2_26 (.CI(n12094), .I0(state_timeout_counter[24]), 
            .I1(VCC_net), .CO(n12095));
    SB_CARRY sub_111_add_2_4 (.CI(n12123), .I0(fifo_state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n12124));
    SB_LUT4 sub_69_add_2_25_lut (.I0(n2075), .I1(state_timeout_counter[23]), 
            .I2(VCC_net), .I3(n12093), .O(n14292)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_69_add_2_10 (.CI(n12078), .I0(state_timeout_counter[8]), 
            .I1(VCC_net), .CO(n12079));
    SB_CARRY sub_69_add_2_25 (.CI(n12093), .I0(state_timeout_counter[23]), 
            .I1(VCC_net), .CO(n12094));
    SB_LUT4 sub_111_add_2_3_lut (.I0(GND_net), .I1(fifo_state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n12122), .O(fifo_state_timeout_counter_5__N_125[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_111_add_2_3 (.CI(n12122), .I0(fifo_state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n12123));
    SB_LUT4 sub_69_add_2_24_lut (.I0(n2075), .I1(state_timeout_counter[22]), 
            .I2(VCC_net), .I3(n12092), .O(n14291)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_111_add_2_2_lut (.I0(GND_net), .I1(fifo_state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(fifo_state_timeout_counter_5__N_125[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_111_add_2_2 (.CI(VCC_net), .I0(fifo_state_timeout_counter[0]), 
            .I1(GND_net), .CO(n12122));
    SB_LUT4 sub_69_add_2_9_lut (.I0(GND_net), .I1(state_timeout_counter[7]), 
            .I2(VCC_net), .I3(n12077), .O(n628[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_9 (.CI(n12077), .I0(state_timeout_counter[7]), 
            .I1(VCC_net), .CO(n12078));
    SB_DFF invert_98_i0 (.Q(reset_all), .C(SLM_CLK_c), .D(n12883));   // src/timing_controller.v(160[5] 229[12])
    SB_LUT4 sub_69_add_2_8_lut (.I0(GND_net), .I1(state_timeout_counter[6]), 
            .I2(VCC_net), .I3(n12076), .O(n628[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR line_of_data_available_91 (.Q(line_of_data_available), .C(SLM_CLK_c), 
            .D(n2), .R(n8043));   // src/timing_controller.v(88[8] 151[4])
    SB_LUT4 i12364_2_lut (.I0(n7), .I1(n8), .I2(GND_net), .I3(GND_net), 
            .O(\aempty_flag_impl.ae_flag_nxt_w ));
    defparam i12364_2_lut.LUT_INIT = 16'h1111;
    SB_DFF invert_98_i4 (.Q(INVERT_c_4), .C(SLM_CLK_c), .D(n1138[4]));   // src/timing_controller.v(160[5] 229[12])
    SB_LUT4 i3430_1_lut (.I0(buffer_switch_done), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4903));   // src/timing_controller.v(160[5] 229[12])
    defparam i3430_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12209_4_lut (.I0(n11566), .I1(fifo_state[2]), .I2(get_next_word), 
            .I3(fifo_state[1]), .O(n14311));
    defparam i12209_4_lut.LUT_INIT = 16'h3011;
    SB_LUT4 i36_3_lut (.I0(n1290), .I1(n11566), .I2(fifo_state[2]), .I3(GND_net), 
            .O(n16));
    defparam i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34_4_lut (.I0(n16), .I1(n14311), .I2(fifo_state[0]), .I3(fifo_state[1]), 
            .O(dc32_fifo_read_enable_N_359));
    defparam i34_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 state_3__I_0_103_Mux_0_i7_4_lut (.I0(state[1]), .I1(n63), .I2(state[2]), 
            .I3(state[0]), .O(n7_adj_1412));   // src/timing_controller.v(160[5] 229[12])
    defparam state_3__I_0_103_Mux_0_i7_4_lut.LUT_INIT = 16'hc535;
    SB_LUT4 state_3__I_0_103_Mux_0_i15_4_lut (.I0(n7_adj_1412), .I1(n9023), 
            .I2(state[3]), .I3(state[0]), .O(state_3__N_83[0]));   // src/timing_controller.v(160[5] 229[12])
    defparam state_3__I_0_103_Mux_0_i15_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i1_2_lut_adj_107 (.I0(fifo_state[2]), .I1(n11566), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_1413));
    defparam i1_2_lut_adj_107.LUT_INIT = 16'h2222;
    SB_LUT4 i12358_4_lut (.I0(fifo_state[1]), .I1(fifo_state_timeout_counter_5__N_125[3]), 
            .I2(fifo_state[0]), .I3(n7_adj_1413), .O(n12868));
    defparam i12358_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i26_3_lut (.I0(n1290), .I1(n11566), .I2(fifo_state[2]), .I3(GND_net), 
            .O(n15));   // src/timing_controller.v(77[11:21])
    defparam i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(fifo_state[0]), .I1(n11540), .I2(fifo_state[1]), 
            .I3(n15), .O(n8321));
    defparam i1_4_lut.LUT_INIT = 16'hcdcc;
    SB_LUT4 i10878_3_lut (.I0(dc32_fifo_almost_empty), .I1(state[3]), .I2(n4688), 
            .I3(GND_net), .O(n1290));
    defparam i10878_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i37_3_lut (.I0(dc32_fifo_full), .I1(get_next_word), .I2(fifo_state[0]), 
            .I3(GND_net), .O(n18));
    defparam i37_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50_3_lut (.I0(n1290), .I1(n11566), .I2(fifo_state[0]), .I3(GND_net), 
            .O(n12988));
    defparam i50_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10934_4_lut (.I0(fifo_state[2]), .I1(n12988), .I2(n18), .I3(fifo_state[1]), 
            .O(n13044));
    defparam i10934_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_4_lut_adj_108 (.I0(fifo_state[2]), .I1(fifo_state[0]), .I2(fifo_state[1]), 
            .I3(n11566), .O(fifo_state_2__N_80[0]));
    defparam i1_4_lut_adj_108.LUT_INIT = 16'h9399;
    SB_LUT4 i1_2_lut_adj_109 (.I0(fifo_state[0]), .I1(n11566), .I2(GND_net), 
            .I3(GND_net), .O(n70));   // src/timing_controller.v(77[11:21])
    defparam i1_2_lut_adj_109.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_110 (.I0(fifo_state[1]), .I1(n11540), .I2(fifo_state[2]), 
            .I3(n70), .O(sc32_fifo_read_enable_N_367));
    defparam i1_4_lut_adj_110.LUT_INIT = 16'hccdc;
    SB_LUT4 i3_4_lut (.I0(fifo_state_timeout_counter[5]), .I1(fifo_state_timeout_counter[1]), 
            .I2(fifo_state_timeout_counter[4]), .I3(fifo_state_timeout_counter[2]), 
            .O(n96));   // src/timing_controller.v(79[11:37])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(n96), .I1(fifo_state_timeout_counter[0]), .I2(fifo_state_timeout_counter[3]), 
            .I3(GND_net), .O(n11566));
    defparam i2_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i12260_2_lut (.I0(get_next_word), .I1(fifo_state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n14276));
    defparam i12260_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_111 (.I0(fifo_state[1]), .I1(n11566), .I2(GND_net), 
            .I3(GND_net), .O(n11));
    defparam i1_2_lut_adj_111.LUT_INIT = 16'heeee;
    SB_CARRY sub_69_add_2_24 (.CI(n12092), .I0(state_timeout_counter[22]), 
            .I1(VCC_net), .CO(n12093));
    SB_LUT4 i20_4_lut (.I0(n11), .I1(n14276), .I2(fifo_state[0]), .I3(fifo_state[2]), 
            .O(sc32_fifo_write_enable_N_366));
    defparam i20_4_lut.LUT_INIT = 16'h05c0;
    SB_LUT4 sub_69_add_2_23_lut (.I0(GND_net), .I1(state_timeout_counter[21]), 
            .I2(VCC_net), .I3(n12091), .O(n628[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_23 (.CI(n12091), .I0(state_timeout_counter[21]), 
            .I1(VCC_net), .CO(n12092));
    SB_CARRY sub_69_add_2_8 (.CI(n12076), .I0(state_timeout_counter[6]), 
            .I1(VCC_net), .CO(n12077));
    SB_LUT4 sub_69_add_2_7_lut (.I0(n4), .I1(state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n12075), .O(n14279)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i12345_2_lut (.I0(state[3]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // src/timing_controller.v(154[8] 230[4])
    defparam i12345_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 sub_69_add_2_22_lut (.I0(n2075), .I1(state_timeout_counter[20]), 
            .I2(VCC_net), .I3(n12090), .O(n14290)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1124_4_lut (.I0(state[3]), .I1(n2334), .I2(n9013), .I3(state[2]), 
            .O(n2252));   // src/timing_controller.v(154[8] 230[4])
    defparam i1124_4_lut.LUT_INIT = 16'h0544;
    SB_CARRY sub_69_add_2_22 (.CI(n12090), .I0(state_timeout_counter[20]), 
            .I1(VCC_net), .CO(n12091));
    SB_LUT4 i6_2_lut (.I0(state_timeout_counter[19]), .I1(state_timeout_counter[21]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // src/timing_controller.v(154[8] 230[4])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut_adj_112 (.I0(state_timeout_counter[22]), .I1(state_timeout_counter[26]), 
            .I2(state_timeout_counter[25]), .I3(state_timeout_counter[28]), 
            .O(n52));   // src/timing_controller.v(154[8] 230[4])
    defparam i20_4_lut_adj_112.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(state_timeout_counter[4]), .I1(state_timeout_counter[16]), 
            .I2(state_timeout_counter[8]), .I3(state_timeout_counter[0]), 
            .O(n56));   // src/timing_controller.v(154[8] 230[4])
    defparam i24_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i22_4_lut (.I0(state_timeout_counter[10]), .I1(state_timeout_counter[17]), 
            .I2(state_timeout_counter[12]), .I3(state_timeout_counter[18]), 
            .O(n54));   // src/timing_controller.v(154[8] 230[4])
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(state_timeout_counter[20]), .I1(state_timeout_counter[1]), 
            .I2(state_timeout_counter[24]), .I3(state_timeout_counter[2]), 
            .O(n55));   // src/timing_controller.v(154[8] 230[4])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(state_timeout_counter[3]), .I1(state_timeout_counter[6]), 
            .I2(state_timeout_counter[5]), .I3(state_timeout_counter[9]), 
            .O(n53));   // src/timing_controller.v(154[8] 230[4])
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(state_timeout_counter[29]), .I1(state_timeout_counter[7]), 
            .I2(state_timeout_counter[30]), .I3(state_timeout_counter[11]), 
            .O(n50));   // src/timing_controller.v(154[8] 230[4])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(state_timeout_counter[13]), .I1(n52), .I2(n38), 
            .I3(state_timeout_counter[14]), .O(n58));   // src/timing_controller.v(154[8] 230[4])
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30_4_lut (.I0(n53), .I1(n55), .I2(n54), .I3(n56), .O(n62));   // src/timing_controller.v(154[8] 230[4])
    defparam i30_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(state_timeout_counter[31]), .I1(state_timeout_counter[23]), 
            .I2(state_timeout_counter[15]), .I3(state_timeout_counter[27]), 
            .O(n49));   // src/timing_controller.v(154[8] 230[4])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31_4_lut (.I0(n49), .I1(n62), .I2(n58), .I3(n50), .O(n63));   // src/timing_controller.v(154[8] 230[4])
    defparam i31_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF invert_98_i1 (.Q(reset_per_frame), .C(SLM_CLK_c), .D(n12884));   // src/timing_controller.v(160[5] 229[12])
    SB_LUT4 i12370_2_lut (.I0(state[3]), .I1(n4688), .I2(GND_net), .I3(GND_net), 
            .O(n4838));
    defparam i12370_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 mux_1055_i1_3_lut (.I0(n14248), .I1(state[1]), .I2(n2180), 
            .I3(GND_net), .O(n2181[0]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1055_i1_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1063_i1_4_lut (.I0(n2181[0]), .I1(state[1]), .I2(n2252), 
            .I3(n12902), .O(n2253[0]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1063_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_DFFESR invert_98_i3 (.Q(UPDATE_c_3), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n14398), .R(n5));   // src/timing_controller.v(160[5] 229[12])
    SB_LUT4 state_3__I_0_103_Mux_1_i15_4_lut_4_lut (.I0(state[0]), .I1(state[1]), 
            .I2(state[3]), .I3(n12914), .O(state_3__N_83[1]));   // src/timing_controller.v(160[5] 229[12])
    defparam state_3__I_0_103_Mux_1_i15_4_lut_4_lut.LUT_INIT = 16'hc6f6;
    SB_LUT4 sub_69_add_2_21_lut (.I0(n2075), .I1(state_timeout_counter[19]), 
            .I2(VCC_net), .I3(n12089), .O(n14289)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_69_add_2_7 (.CI(n12075), .I0(state_timeout_counter[5]), 
            .I1(VCC_net), .CO(n12076));
    SB_LUT4 i1_2_lut_adj_113 (.I0(fifo_state[2]), .I1(n1290), .I2(GND_net), 
            .I3(GND_net), .O(n17));
    defparam i1_2_lut_adj_113.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_114 (.I0(fifo_state[0]), .I1(fifo_state[1]), .I2(n17), 
            .I3(n12900), .O(n8325));
    defparam i1_4_lut_adj_114.LUT_INIT = 16'hba32;
    SB_LUT4 i1_2_lut_adj_115 (.I0(fifo_state[1]), .I1(n12865), .I2(GND_net), 
            .I3(GND_net), .O(n12866));   // src/timing_controller.v(88[8] 151[4])
    defparam i1_2_lut_adj_115.LUT_INIT = 16'h4444;
    SB_LUT4 i123_4_lut (.I0(fifo_state[2]), .I1(fifo_state[0]), .I2(fifo_state_timeout_counter[0]), 
            .I3(n4_adj_1414), .O(n94));   // src/timing_controller.v(77[11:21])
    defparam i123_4_lut.LUT_INIT = 16'heece;
    SB_LUT4 i1_2_lut_adj_116 (.I0(n96), .I1(fifo_state_timeout_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1414));   // src/timing_controller.v(79[11:37])
    defparam i1_2_lut_adj_116.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_4_lut (.I0(fifo_state[1]), .I1(fifo_state[0]), .I2(fifo_state[2]), 
            .I3(get_next_word), .O(n11540));   // src/timing_controller.v(88[8] 151[4])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i25_1_lut (.I0(dc32_fifo_read_enable), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // src/top.v(482[26:47])
    defparam i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[3]), .I1(n63), .I2(state[1]), .I3(state[2]), 
            .O(n12908));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_adj_117 (.I0(state[0]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n12882));
    defparam i1_2_lut_adj_117.LUT_INIT = 16'h2222;
    SB_LUT4 i7296_2_lut (.I0(dc32_fifo_full), .I1(fifo_state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // src/timing_controller.v(93[5] 150[12])
    defparam i7296_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_118 (.I0(fifo_state[2]), .I1(fifo_state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n8043));   // src/timing_controller.v(88[8] 151[4])
    defparam i1_2_lut_adj_118.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_119 (.I0(state[1]), .I1(state[3]), 
            .I2(state[0]), .I3(state[2]), .O(n12883));   // src/timing_controller.v(160[5] 229[12])
    defparam i1_2_lut_3_lut_4_lut_adj_119.LUT_INIT = 16'h0010;
    SB_LUT4 i3945_2_lut_3_lut (.I0(state[3]), .I1(n4688), .I2(n2252), 
            .I3(GND_net), .O(n5419));   // src/timing_controller.v(154[8] 230[4])
    defparam i3945_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i12342_3_lut_4_lut (.I0(state[3]), .I1(n4688), .I2(n2252), 
            .I3(n4), .O(n5404));
    defparam i12342_3_lut_4_lut.LUT_INIT = 16'h7077;
    SB_LUT4 i12287_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n14398));   // src/timing_controller.v(160[5] 229[12])
    defparam i12287_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_120 (.I0(state[0]), .I1(n63), .I2(state[3]), 
            .I3(state[2]), .O(n12902));   // src/timing_controller.v(154[8] 230[4])
    defparam i1_2_lut_3_lut_4_lut_adj_120.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_3_lut_adj_121 (.I0(n9015), .I1(state[3]), .I2(n63), 
            .I3(GND_net), .O(n4936));
    defparam i1_2_lut_3_lut_adj_121.LUT_INIT = 16'hdfdf;
    SB_LUT4 i1_2_lut_adj_122 (.I0(fifo_state[2]), .I1(get_next_word), .I2(GND_net), 
            .I3(GND_net), .O(n12900));   // src/timing_controller.v(88[8] 151[4])
    defparam i1_2_lut_adj_122.LUT_INIT = 16'h4444;
>>>>>>> Stashed changes
    
endmodule
//
// Verilog Description of module bluejay_data
//

<<<<<<< Updated upstream
module timing_controller (state, SLM_CLK_c, n1879, GND_net, n10514, 
            VCC_net, n10808, reset_per_frame, n1774, n7386, INVERT_c_3, 
            buffer_switch_done, n4245, n7568, n7590, n4192, n63, 
            n10831, UPDATE_c_2) /* synthesis syn_module_defined=1 */ ;
    output [3:0]state;
=======
module bluejay_data (VCC_net, DEBUG_6_c, SLM_CLK_c, GND_net, n4903, 
            buffer_switch_done, n6968, DEBUG_8_c, buffer_switch_done_latched, 
            n934, n12261, n1013, bluejay_data_out_31__N_920, bluejay_data_out_31__N_921, 
            bluejay_data_out_31__N_922, SYNC_c, DATA10_c_10, n5367, 
            line_of_data_available, DATA9_c_9, n5366, DATA11_c_11, n5365, 
            DATA12_c_12, n5364, DATA13_c_13, n5363, DATA14_c_14, n5362, 
            DATA8_c_8, n5361, DATA15_c_15, n5360, DATA16_c_16, n5359, 
            DATA7_c_7, n5358, DATA17_c_17, n5357, DATA18_c_18, n5356, 
            DATA6_c_6, n5355, DATA19_c_19, n5354, DATA20_c_20, n5353, 
            DATA5_c_5, n5352, DATA21_c_21, n5351, DATA22_c_22, n5350, 
            DATA4_c_4, n5349, DATA23_c_23, n5348, DATA24_c_24, n5347, 
            DATA3_c_3, n5346, DATA25_c_25, n5345, DATA26_c_26, n5344, 
            DATA2_c_2, n5343, DATA27_c_27, n5342, n5573, get_next_word, 
            DATA28_c_28, n5341, DATA1_c_1, n5340, DATA29_c_29, n5339, 
            DATA30_c_30, n5338, DATA31_c_31, n5337, sc32_fifo_almost_empty) /* synthesis syn_module_defined=1 */ ;
    input VCC_net;
    output DEBUG_6_c;
>>>>>>> Stashed changes
    input SLM_CLK_c;
    input n1879;
    input GND_net;
<<<<<<< Updated upstream
    input n10514;
    input VCC_net;
    input n10808;
    output reset_per_frame;
    input n1774;
    input n7386;
    output INVERT_c_3;
    output buffer_switch_done;
    output n4245;
    output n7568;
    input n7590;
    output n4192;
    output n63;
    output n10831;
    output UPDATE_c_2;
=======
    input n4903;
    input buffer_switch_done;
    input n6968;
    output DEBUG_8_c;
    input buffer_switch_done_latched;
    output n934;
    input n12261;
    output n1013;
    output bluejay_data_out_31__N_920;
    output bluejay_data_out_31__N_921;
    output bluejay_data_out_31__N_922;
    output SYNC_c;
    output DATA10_c_10;
    input n5367;
    input line_of_data_available;
    output DATA9_c_9;
    input n5366;
    output DATA11_c_11;
    input n5365;
    output DATA12_c_12;
    input n5364;
    output DATA13_c_13;
    input n5363;
    output DATA14_c_14;
    input n5362;
    output DATA8_c_8;
    input n5361;
    output DATA15_c_15;
    input n5360;
    output DATA16_c_16;
    input n5359;
    output DATA7_c_7;
    input n5358;
    output DATA17_c_17;
    input n5357;
    output DATA18_c_18;
    input n5356;
    output DATA6_c_6;
    input n5355;
    output DATA19_c_19;
    input n5354;
    output DATA20_c_20;
    input n5353;
    output DATA5_c_5;
    input n5352;
    output DATA21_c_21;
    input n5351;
    output DATA22_c_22;
    input n5350;
    output DATA4_c_4;
    input n5349;
    output DATA23_c_23;
    input n5348;
    output DATA24_c_24;
    input n5347;
    output DATA3_c_3;
    input n5346;
    output DATA25_c_25;
    input n5345;
    output DATA26_c_26;
    input n5344;
    output DATA2_c_2;
    input n5343;
    output DATA27_c_27;
    input n5342;
    input n5573;
    output get_next_word;
    output DATA28_c_28;
    input n5341;
    output DATA1_c_1;
    input n5340;
    output DATA29_c_29;
    input n5339;
    output DATA30_c_30;
    input n5338;
    output DATA31_c_31;
    input n5337;
    input sc32_fifo_almost_empty;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [8:0]n74;
    
    wire n5, n12904, n8, n12597, n12150;
    wire [10:0]v_counter;   // src/bluejay_data.v(51[12:21])
    
    wire n12151, valid_N_925;
    wire [10:0]v_counter_10__N_900;
    
    wire n12149, n12405;
    wire [7:0]state_timeout_counter;   // src/bluejay_data.v(52[11:32])
    
    wire n5516, n12429, n5515, n12834, n5514, n12485, n5513, n5_adj_1403, 
        n12453, n9, n5511, n12563, n5388, n12148;
    wire [15:0]n998;
    
    wire n5007, n12147, n3, n7, n7_adj_1404;
    wire [3:0]n99;
    
    wire n8_adj_1405, n12064, n12065, n12146, n12145, n12144, n12061, 
        n12059, n12060, n12062, n12063, n32, n3_adj_1406, n6, 
        n1537, n1307, n12842, n1052, bluejay_data_out_31__N_919, n3477, 
        n3479, n1061, n3481, n1065, n3483, n3_adj_1407, n4, n6_adj_1408, 
        n12837, n4_adj_1409, n12817, n12916, n4_adj_1410, n12823, 
        n12905, n12153, n12152, n13014, n4_adj_1411, n12239, n68;
    
    SB_LUT4 i2_4_lut (.I0(n74[0]), .I1(n5), .I2(n12904), .I3(n8), .O(n12597));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2_4_lut.LUT_INIT = 16'hffec;
    SB_CARRY sub_123_add_2_9 (.CI(n12150), .I0(v_counter[7]), .I1(VCC_net), 
            .CO(n12151));
    SB_DFFN valid_66 (.Q(DEBUG_6_c), .C(SLM_CLK_c), .D(valid_N_925));   // src/bluejay_data.v(134[8] 156[4])
    SB_LUT4 sub_123_add_2_8_lut (.I0(GND_net), .I1(v_counter[6]), .I2(VCC_net), 
            .I3(n12149), .O(v_counter_10__N_900[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_123_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS state_timeout_counter_i0_i7 (.Q(state_timeout_counter[7]), .C(SLM_CLK_c), 
            .E(n4903), .D(n12405), .S(n5516));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS state_timeout_counter_i0_i6 (.Q(state_timeout_counter[6]), .C(SLM_CLK_c), 
            .E(n4903), .D(n12429), .S(n5515));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS state_timeout_counter_i0_i5 (.Q(state_timeout_counter[5]), .C(SLM_CLK_c), 
            .E(n4903), .D(n12834), .S(n5514));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(SLM_CLK_c), 
            .E(n4903), .D(n12485), .S(n5513));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(SLM_CLK_c), 
            .E(n4903), .D(n5_adj_1403), .S(n12453));   // src/bluejay_data.v(56[8] 131[4])
    SB_CARRY sub_123_add_2_8 (.CI(n12149), .I0(v_counter[6]), .I1(VCC_net), 
            .CO(n12150));
    SB_DFFESS state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(SLM_CLK_c), 
            .E(n4903), .D(n9), .S(n5511));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(SLM_CLK_c), 
            .E(n4903), .D(n12563), .S(n5388));   // src/bluejay_data.v(56[8] 131[4])
    SB_LUT4 sub_123_add_2_7_lut (.I0(GND_net), .I1(v_counter[5]), .I2(VCC_net), 
            .I3(n12148), .O(v_counter_10__N_900[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_123_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_123_add_2_7 (.CI(n12148), .I0(v_counter[5]), .I1(VCC_net), 
            .CO(n12149));
    SB_LUT4 i1_2_lut (.I0(n998[9]), .I1(buffer_switch_done), .I2(GND_net), 
            .I3(GND_net), .O(n5007));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 sub_123_add_2_6_lut (.I0(GND_net), .I1(v_counter[4]), .I2(VCC_net), 
            .I3(n12147), .O(v_counter_10__N_900[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_123_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFN bluejay_data_out_i1 (.Q(DEBUG_8_c), .C(SLM_CLK_c), .D(n6968));   // src/bluejay_data.v(134[8] 156[4])
    SB_LUT4 i1_2_lut_3_lut (.I0(n998[2]), .I1(buffer_switch_done_latched), 
            .I2(state_timeout_counter[0]), .I3(GND_net), .O(n5));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1_2_lut_3_lut_adj_79 (.I0(n998[2]), .I1(buffer_switch_done_latched), 
            .I2(state_timeout_counter[1]), .I3(GND_net), .O(n3));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_3_lut_adj_79.LUT_INIT = 16'h2020;
    SB_LUT4 i1_2_lut_3_lut_adj_80 (.I0(n998[2]), .I1(buffer_switch_done_latched), 
            .I2(state_timeout_counter[7]), .I3(GND_net), .O(n7));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_3_lut_adj_80.LUT_INIT = 16'h2020;
    SB_LUT4 i1_2_lut_3_lut_adj_81 (.I0(n998[2]), .I1(buffer_switch_done_latched), 
            .I2(state_timeout_counter[4]), .I3(GND_net), .O(n7_adj_1404));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_3_lut_adj_81.LUT_INIT = 16'h2020;
    SB_LUT4 i1_3_lut_4_lut (.I0(n99[2]), .I1(n934), .I2(n74[0]), .I3(n998[9]), 
            .O(n8));   // src/bluejay_data.v(107[17] 116[20])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 i1_3_lut_4_lut_adj_82 (.I0(n99[2]), .I1(n934), .I2(n74[1]), 
            .I3(n998[9]), .O(n8_adj_1405));   // src/bluejay_data.v(107[17] 116[20])
    defparam i1_3_lut_4_lut_adj_82.LUT_INIT = 16'hf200;
    SB_CARRY sub_121_add_2_8 (.CI(n12064), .I0(state_timeout_counter[6]), 
            .I1(VCC_net), .CO(n12065));
    SB_CARRY sub_123_add_2_6 (.CI(n12147), .I0(v_counter[4]), .I1(VCC_net), 
            .CO(n12148));
    SB_LUT4 sub_123_add_2_5_lut (.I0(GND_net), .I1(v_counter[3]), .I2(VCC_net), 
            .I3(n12146), .O(v_counter_10__N_900[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_123_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_123_add_2_5 (.CI(n12146), .I0(v_counter[3]), .I1(VCC_net), 
            .CO(n12147));
    SB_LUT4 sub_123_add_2_4_lut (.I0(GND_net), .I1(v_counter[2]), .I2(VCC_net), 
            .I3(n12145), .O(v_counter_10__N_900[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_123_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_123_add_2_4 (.CI(n12145), .I0(v_counter[2]), .I1(VCC_net), 
            .CO(n12146));
    SB_LUT4 sub_123_add_2_3_lut (.I0(GND_net), .I1(v_counter[1]), .I2(VCC_net), 
            .I3(n12144), .O(v_counter_10__N_900[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_123_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_121_add_2_5_lut (.I0(GND_net), .I1(state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n12061), .O(n74[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_121_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_123_add_2_3 (.CI(n12144), .I0(v_counter[1]), .I1(VCC_net), 
            .CO(n12145));
    SB_LUT4 sub_123_add_2_2_lut (.I0(GND_net), .I1(v_counter[0]), .I2(n934), 
            .I3(VCC_net), .O(v_counter_10__N_900[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_123_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR v_counter_i10 (.Q(v_counter[10]), .C(SLM_CLK_c), .E(n5007), 
            .D(v_counter_10__N_900[10]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_LUT4 sub_121_add_2_3_lut (.I0(GND_net), .I1(state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n12059), .O(n74[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_121_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR v_counter_i9 (.Q(v_counter[9]), .C(SLM_CLK_c), .E(n5007), 
            .D(v_counter_10__N_900[9]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i8 (.Q(v_counter[8]), .C(SLM_CLK_c), .E(n5007), 
            .D(v_counter_10__N_900[8]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i7 (.Q(v_counter[7]), .C(SLM_CLK_c), .E(n5007), 
            .D(v_counter_10__N_900[7]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i6 (.Q(v_counter[6]), .C(SLM_CLK_c), .E(n5007), 
            .D(v_counter_10__N_900[6]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_CARRY sub_123_add_2_2 (.CI(VCC_net), .I0(v_counter[0]), .I1(n934), 
            .CO(n12144));
    SB_DFFESS v_counter_i5 (.Q(v_counter[5]), .C(SLM_CLK_c), .E(n5007), 
            .D(v_counter_10__N_900[5]), .S(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i4 (.Q(v_counter[4]), .C(SLM_CLK_c), .E(n5007), 
            .D(v_counter_10__N_900[4]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i3 (.Q(v_counter[3]), .C(SLM_CLK_c), .E(n5007), 
            .D(v_counter_10__N_900[3]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i2 (.Q(v_counter[2]), .C(SLM_CLK_c), .E(n5007), 
            .D(v_counter_10__N_900[2]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i1 (.Q(v_counter[1]), .C(SLM_CLK_c), .E(n5007), 
            .D(v_counter_10__N_900[1]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_CARRY sub_121_add_2_3 (.CI(n12059), .I0(state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n12060));
    SB_DFFESS state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(SLM_CLK_c), 
            .E(n4903), .D(n12597), .S(n5388));   // src/bluejay_data.v(56[8] 131[4])
    SB_CARRY sub_121_add_2_5 (.CI(n12061), .I0(state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n12062));
    SB_LUT4 sub_121_add_2_2_lut (.I0(GND_net), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n74[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_121_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_121_add_2_4_lut (.I0(GND_net), .I1(state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n12060), .O(n74[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_121_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_121_add_2_2 (.CI(VCC_net), .I0(state_timeout_counter[0]), 
            .I1(GND_net), .CO(n12059));
    SB_CARRY sub_121_add_2_4 (.CI(n12060), .I0(state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n12061));
    SB_DFFESR v_counter_i0 (.Q(v_counter[0]), .C(SLM_CLK_c), .E(n5007), 
            .D(v_counter_10__N_900[0]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_LUT4 i2_4_lut_adj_83 (.I0(n74[1]), .I1(n3), .I2(n12904), .I3(n8_adj_1405), 
            .O(n12563));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2_4_lut_adj_83.LUT_INIT = 16'hffec;
    SB_CARRY sub_121_add_2_6 (.CI(n12062), .I0(state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n12063));
    SB_LUT4 i1_2_lut_adj_84 (.I0(n998[2]), .I1(state_timeout_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_84.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_85 (.I0(buffer_switch_done_latched), .I1(n74[2]), 
            .I2(n32), .I3(n3_adj_1406), .O(n6));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2_4_lut_adj_85.LUT_INIT = 16'hfefa;
    SB_LUT4 i3_4_lut (.I0(n74[2]), .I1(n1537), .I2(n998[5]), .I3(n1307), 
            .O(n9));   // src/bluejay_data.v(66[9] 129[16])
    defparam i3_4_lut.LUT_INIT = 16'ha8f8;
    SB_DFFSR state_FSM_i2 (.Q(n1013), .C(SLM_CLK_c), .D(n12261), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i3 (.Q(n998[2]), .C(SLM_CLK_c), .D(n12842), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i4 (.Q(bluejay_data_out_31__N_919), .C(SLM_CLK_c), 
            .D(n1052), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i5 (.Q(n998[4]), .C(SLM_CLK_c), .D(n3477), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i6 (.Q(n998[5]), .C(SLM_CLK_c), .D(n3479), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i7 (.Q(bluejay_data_out_31__N_920), .C(SLM_CLK_c), 
            .D(n1061), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i8 (.Q(bluejay_data_out_31__N_921), .C(SLM_CLK_c), 
            .D(n3481), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i9 (.Q(bluejay_data_out_31__N_922), .C(SLM_CLK_c), 
            .D(n1065), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i10 (.Q(n998[9]), .C(SLM_CLK_c), .D(n3483), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFN sync_68 (.Q(SYNC_c), .C(SLM_CLK_c), .D(bluejay_data_out_31__N_919));   // src/bluejay_data.v(134[8] 156[4])
    SB_LUT4 i2_3_lut (.I0(n998[2]), .I1(buffer_switch_done_latched), .I2(state_timeout_counter[3]), 
            .I3(GND_net), .O(n3_adj_1407));   // src/bluejay_data.v(56[8] 131[4])
    defparam i2_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1_4_lut (.I0(n4903), .I1(n1537), .I2(n3_adj_1407), .I3(n74[3]), 
            .O(n12453));   // src/bluejay_data.v(56[8] 131[4])
    defparam i1_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_2_lut_adj_86 (.I0(n74[3]), .I1(n4), .I2(GND_net), .I3(GND_net), 
            .O(n5_adj_1403));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_86.LUT_INIT = 16'h8888;
    SB_LUT4 i4039_4_lut (.I0(n4903), .I1(n74[4]), .I2(n7_adj_1404), .I3(n1537), 
            .O(n5513));   // src/bluejay_data.v(56[8] 131[4])
    defparam i4039_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_2_lut_adj_87 (.I0(n74[4]), .I1(n4), .I2(GND_net), .I3(GND_net), 
            .O(n12485));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_87.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_88 (.I0(buffer_switch_done_latched), .I1(n998[2]), 
            .I2(n6_adj_1408), .I3(state_timeout_counter[5]), .O(n12834));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_4_lut_adj_88.LUT_INIT = 16'hfefa;
    SB_DFFNESR bluejay_data_out_i11 (.Q(DATA10_c_10), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5367));   // src/bluejay_data.v(134[8] 156[4])
    SB_LUT4 i1_4_lut_adj_89 (.I0(n74[6]), .I1(n998[2]), .I2(n1537), .I3(state_timeout_counter[6]), 
            .O(n12837));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_4_lut_adj_89.LUT_INIT = 16'heca0;
    SB_LUT4 i1_2_lut_adj_90 (.I0(n74[6]), .I1(n4), .I2(GND_net), .I3(GND_net), 
            .O(n12429));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_90.LUT_INIT = 16'h8888;
    SB_LUT4 i548_2_lut (.I0(line_of_data_available), .I1(n934), .I2(GND_net), 
            .I3(GND_net), .O(n1307));   // src/bluejay_data.v(120[17] 127[20])
    defparam i548_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_91 (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[7]), 
            .I2(state_timeout_counter[2]), .I3(state_timeout_counter[6]), 
            .O(n4_adj_1409));   // src/bluejay_data.v(107[21:49])
    defparam i1_4_lut_adj_91.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_92 (.I0(state_timeout_counter[4]), .I1(n4_adj_1409), 
            .I2(state_timeout_counter[3]), .I3(GND_net), .O(n12817));   // src/bluejay_data.v(107[21:49])
    defparam i2_3_lut_adj_92.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_93 (.I0(v_counter[5]), .I1(v_counter[8]), .I2(v_counter[2]), 
            .I3(v_counter[4]), .O(n12916));
    defparam i3_4_lut_adj_93.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_94 (.I0(v_counter[3]), .I1(v_counter[0]), .I2(v_counter[6]), 
            .I3(v_counter[1]), .O(n4_adj_1410));   // src/bluejay_data.v(109[25:41])
    defparam i1_4_lut_adj_94.LUT_INIT = 16'hfffb;
    SB_LUT4 i2_4_lut_adj_95 (.I0(v_counter[10]), .I1(n4_adj_1410), .I2(v_counter[7]), 
            .I3(v_counter[9]), .O(n12823));   // src/bluejay_data.v(109[25:41])
    defparam i2_4_lut_adj_95.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_96 (.I0(state_timeout_counter[5]), .I1(state_timeout_counter[0]), 
            .I2(n12817), .I3(GND_net), .O(n934));   // src/bluejay_data.v(107[21:49])
    defparam i2_3_lut_adj_96.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_adj_97 (.I0(n12823), .I1(n12916), .I2(GND_net), .I3(GND_net), 
            .O(n99[2]));   // src/bluejay_data.v(109[25:41])
    defparam i1_2_lut_adj_97.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_98 (.I0(bluejay_data_out_31__N_921), .I1(n998[4]), 
            .I2(n1013), .I3(GND_net), .O(n1537));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2_3_lut_adj_98.LUT_INIT = 16'hfefe;
    SB_LUT4 i4042_4_lut (.I0(n4903), .I1(n74[7]), .I2(n7), .I3(n1537), 
            .O(n5516));   // src/bluejay_data.v(56[8] 131[4])
    defparam i4042_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_2_lut_adj_99 (.I0(n74[7]), .I1(n4), .I2(GND_net), .I3(GND_net), 
            .O(n12405));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_99.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_100 (.I0(bluejay_data_out_31__N_921), .I1(bluejay_data_out_31__N_922), 
            .I2(GND_net), .I3(GND_net), .O(valid_N_925));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_100.LUT_INIT = 16'heeee;
    SB_DFFNESR bluejay_data_out_i10 (.Q(DATA9_c_9), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5366));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i12 (.Q(DATA11_c_11), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5365));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i13 (.Q(DATA12_c_12), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5364));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i14 (.Q(DATA13_c_13), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5363));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i15 (.Q(DATA14_c_14), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5362));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i9 (.Q(DATA8_c_8), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5361));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i16 (.Q(DATA15_c_15), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5360));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i17 (.Q(DATA16_c_16), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5359));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i8 (.Q(DATA7_c_7), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5358));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i18 (.Q(DATA17_c_17), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5357));   // src/bluejay_data.v(134[8] 156[4])
    SB_LUT4 sub_121_add_2_7_lut (.I0(n12905), .I1(state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n12063), .O(n6_adj_1408)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_121_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_DFFNESR bluejay_data_out_i19 (.Q(DATA18_c_18), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5356));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i7 (.Q(DATA6_c_6), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5355));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i20 (.Q(DATA19_c_19), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5354));   // src/bluejay_data.v(134[8] 156[4])
    SB_LUT4 sub_123_add_2_12_lut (.I0(GND_net), .I1(v_counter[10]), .I2(VCC_net), 
            .I3(n12153), .O(v_counter_10__N_900[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_123_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_121_add_2_9_lut (.I0(GND_net), .I1(state_timeout_counter[7]), 
            .I2(VCC_net), .I3(n12065), .O(n74[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_121_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_121_add_2_8_lut (.I0(GND_net), .I1(state_timeout_counter[6]), 
            .I2(VCC_net), .I3(n12064), .O(n74[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_121_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_123_add_2_11_lut (.I0(GND_net), .I1(v_counter[9]), .I2(VCC_net), 
            .I3(n12152), .O(v_counter_10__N_900[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_123_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_123_add_2_11 (.CI(n12152), .I0(v_counter[9]), .I1(VCC_net), 
            .CO(n12153));
    SB_LUT4 sub_121_add_2_6_lut (.I0(GND_net), .I1(state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n12062), .O(n74[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_121_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_123_add_2_10_lut (.I0(GND_net), .I1(v_counter[8]), .I2(VCC_net), 
            .I3(n12151), .O(v_counter_10__N_900[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_123_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_DFFNESR bluejay_data_out_i21 (.Q(DATA20_c_20), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5353));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i6 (.Q(DATA5_c_5), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5352));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i22 (.Q(DATA21_c_21), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5351));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i23 (.Q(DATA22_c_22), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5350));   // src/bluejay_data.v(134[8] 156[4])
    SB_CARRY sub_121_add_2_7 (.CI(n12063), .I0(state_timeout_counter[5]), 
            .I1(VCC_net), .CO(n12064));
    SB_DFFNESR bluejay_data_out_i5 (.Q(DATA4_c_4), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5349));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i24 (.Q(DATA23_c_23), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5348));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i25 (.Q(DATA24_c_24), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5347));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i4 (.Q(DATA3_c_3), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5346));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i26 (.Q(DATA25_c_25), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5345));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i27 (.Q(DATA26_c_26), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5344));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i3 (.Q(DATA2_c_2), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5343));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i28 (.Q(DATA27_c_27), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5342));   // src/bluejay_data.v(134[8] 156[4])
    SB_LUT4 i2024_3_lut_4_lut (.I0(buffer_switch_done_latched), .I1(n934), 
            .I2(bluejay_data_out_31__N_919), .I3(n998[4]), .O(n3477));   // src/bluejay_data.v(62[9] 65[12])
    defparam i2024_3_lut_4_lut.LUT_INIT = 16'hf4f0;
    SB_LUT4 i1_3_lut_4_lut_adj_101 (.I0(buffer_switch_done_latched), .I1(n934), 
            .I2(bluejay_data_out_31__N_922), .I3(n998[9]), .O(n3483));   // src/bluejay_data.v(62[9] 65[12])
    defparam i1_3_lut_4_lut_adj_101.LUT_INIT = 16'hf4f0;
    SB_LUT4 reduce_or_361_i1_4_lut_4_lut (.I0(n934), .I1(line_of_data_available), 
            .I2(n998[4]), .I3(n998[5]), .O(n1061));   // src/bluejay_data.v(69[17] 76[20])
    defparam reduce_or_361_i1_4_lut_4_lut.LUT_INIT = 16'h5450;
    SB_LUT4 i353_2_lut_3_lut (.I0(n934), .I1(line_of_data_available), .I2(n1013), 
            .I3(GND_net), .O(n1052));   // src/bluejay_data.v(69[17] 76[20])
    defparam i353_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_DFFN get_next_word_67 (.Q(get_next_word), .C(SLM_CLK_c), .D(n5573));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i29 (.Q(DATA28_c_28), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5341));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i2 (.Q(DATA1_c_1), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5340));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i30 (.Q(DATA29_c_29), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5339));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i31 (.Q(DATA30_c_30), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5338));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i32 (.Q(DATA31_c_31), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5337));   // src/bluejay_data.v(134[8] 156[4])
    SB_CARRY sub_123_add_2_10 (.CI(n12151), .I0(v_counter[8]), .I1(VCC_net), 
            .CO(n12152));
    SB_LUT4 sub_123_add_2_9_lut (.I0(GND_net), .I1(v_counter[7]), .I2(VCC_net), 
            .I3(n12150), .O(v_counter_10__N_900[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_123_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i366_2_lut_3_lut (.I0(n934), .I1(sc32_fifo_almost_empty), .I2(bluejay_data_out_31__N_921), 
            .I3(GND_net), .O(n1065));   // src/bluejay_data.v(66[9] 129[16])
    defparam i366_2_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 i4041_3_lut_3_lut (.I0(buffer_switch_done), .I1(buffer_switch_done_latched), 
            .I2(n12837), .I3(GND_net), .O(n5515));   // src/bluejay_data.v(56[8] 131[4])
    defparam i4041_3_lut_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i4040_2_lut_2_lut (.I0(buffer_switch_done), .I1(bluejay_data_out_31__N_920), 
            .I2(GND_net), .I3(GND_net), .O(n5514));   // src/bluejay_data.v(56[8] 131[4])
    defparam i4040_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4037_4_lut_4_lut (.I0(buffer_switch_done), .I1(bluejay_data_out_31__N_922), 
            .I2(n6), .I3(bluejay_data_out_31__N_920), .O(n5511));   // src/bluejay_data.v(56[8] 131[4])
    defparam i4037_4_lut_4_lut.LUT_INIT = 16'h5554;
    SB_LUT4 i3914_3_lut_3_lut (.I0(buffer_switch_done), .I1(bluejay_data_out_31__N_920), 
            .I2(bluejay_data_out_31__N_919), .I3(GND_net), .O(n5388));   // src/bluejay_data.v(56[8] 131[4])
    defparam i3914_3_lut_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_4_lut_adj_102 (.I0(n998[2]), .I1(n13014), .I2(n1013), .I3(n1307), 
            .O(n12842));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_4_lut_adj_102.LUT_INIT = 16'hbbfb;
    SB_LUT4 i10905_4_lut (.I0(n12823), .I1(state_timeout_counter[5]), .I2(n4_adj_1411), 
            .I3(n12916), .O(n13014));
    defparam i10905_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(n998[9]), .I1(n12817), .I2(state_timeout_counter[0]), 
            .I3(GND_net), .O(n4_adj_1411));
    defparam i1_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i2026_4_lut (.I0(n12239), .I1(n998[9]), .I2(n99[2]), .I3(n934), 
            .O(n3479));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2026_4_lut.LUT_INIT = 16'haaea;
    SB_LUT4 i2_4_lut_adj_103 (.I0(buffer_switch_done_latched), .I1(n934), 
            .I2(n998[5]), .I3(line_of_data_available), .O(n12239));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2_4_lut_adj_103.LUT_INIT = 16'h4050;
    SB_LUT4 i2028_4_lut (.I0(buffer_switch_done_latched), .I1(bluejay_data_out_31__N_920), 
            .I2(n68), .I3(bluejay_data_out_31__N_921), .O(n3481));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2028_4_lut.LUT_INIT = 16'hcdcc;
    SB_LUT4 i19_2_lut (.I0(n934), .I1(sc32_fifo_almost_empty), .I2(GND_net), 
            .I3(GND_net), .O(n68));   // src/bluejay_data.v(97[21:87])
    defparam i19_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_104 (.I0(n3_adj_1406), .I1(n12904), .I2(GND_net), 
            .I3(GND_net), .O(n12905));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_104.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n12823), .I1(n12916), .I2(n934), 
            .I3(n998[9]), .O(n3_adj_1406));   // src/bluejay_data.v(107[17] 116[20])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hf100;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_105 (.I0(n998[5]), .I1(line_of_data_available), 
            .I2(n934), .I3(n1537), .O(n12904));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_3_lut_4_lut_adj_105.LUT_INIT = 16'hffa8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_106 (.I0(n998[5]), .I1(line_of_data_available), 
            .I2(n934), .I3(n3_adj_1406), .O(n4));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_3_lut_4_lut_adj_106.LUT_INIT = 16'hffa8;
    
endmodule
//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=20) 
//

module \uart_rx(CLKS_PER_BIT=20)  (SLM_CLK_c, r_Rx_Data, r_Bit_Index, 
            n4790, GND_net, n4, n6967, pc_data_rx, VCC_net, debug_led3, 
            n6956, n6909, n6908, n6907, n6906, n6905, n6904, n6903, 
            n13008, n13034, UART_RX_c, n4787, n4_adj_9, n4_adj_10, 
            n4794) /* synthesis syn_module_defined=1 */ ;
    input SLM_CLK_c;
    output r_Rx_Data;
    output [2:0]r_Bit_Index;
    output n4790;
    input GND_net;
    output n4;
    input n6967;
    output [7:0]pc_data_rx;
    input VCC_net;
    output debug_led3;
    input n6956;
    input n6909;
    input n6908;
    input n6907;
    input n6906;
    input n6905;
    input n6904;
    input n6903;
    output n13008;
    output n13034;
    input UART_RX_c;
    output n4787;
    output n4_adj_9;
    output n4_adj_10;
    output n4794;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [2:0]r_SM_Main;   // src/uart_rx.v(36[17:26])
    wire [2:0]r_SM_Main_2__N_950;
    
    wire n4693, n3, r_Rx_Data_R;
    wire [2:0]r_Bit_Index_c;   // src/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main_2__N_956;
    
    wire n4_adj_1398, n13024, n5532, n6, n4913;
    wire [9:0]n45;
    wire [9:0]r_Clock_Count;   // src/uart_rx.v(32[17:30])
    
    wire n12195, n12194, n12193, n12192;
    wire [2:0]n340;
    
    wire n12411, n9011, n12191, n12190, n12189, n12188, n12187, 
        n12875, n9053, n4691, n8, n6_adj_1399, n4_adj_1400, n9043, 
        n1, n4870;
    
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main_2__N_950[2]), .O(n4693));   // src/uart_rx.v(52[7] 143[14])
    defparam i2_4_lut.LUT_INIT = 16'hfdff;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(SLM_CLK_c), .D(n3), .R(r_SM_Main[2]));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(SLM_CLK_c), .D(r_Rx_Data_R));   // src/uart_rx.v(41[10] 45[8])
    SB_LUT4 i1_2_lut (.I0(r_Bit_Index[0]), .I1(n4693), .I2(GND_net), .I3(GND_net), 
            .O(n4790));   // src/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_150_i4_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // src/uart_rx.v(97[17:39])
    defparam equal_150_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_76 (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_956[0]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1398));
    defparam i1_2_lut_adj_76.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n13024), .I2(r_SM_Main_2__N_950[2]), 
            .I3(r_SM_Main[1]), .O(n5532));
    defparam i1_4_lut.LUT_INIT = 16'h5011;
    SB_LUT4 i2_2_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_956[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12335_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6), 
            .I3(r_SM_Main[0]), .O(n4913));   // src/uart_rx.v(52[7] 143[14])
    defparam i12335_4_lut.LUT_INIT = 16'h4555;
    SB_LUT4 r_Clock_Count_1439_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[9]), .I3(n12195), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1439_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1439_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n12194), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1439_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1439_add_4_10 (.CI(n12194), .I0(GND_net), .I1(r_Clock_Count[8]), 
            .CO(n12195));
    SB_LUT4 r_Clock_Count_1439_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n12193), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1439_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1439_add_4_9 (.CI(n12193), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n12194));
    SB_LUT4 r_Clock_Count_1439_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n12192), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1439_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1600_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n340[1]));   // src/uart_rx.v(102[36:51])
    defparam i1600_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Rx_Byte_i0 (.Q(pc_data_rx[0]), .C(SLM_CLK_c), .D(n6967));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Rx_DV_52 (.Q(debug_led3), .C(SLM_CLK_c), .E(VCC_net), .D(n12411));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n6956));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(pc_data_rx[1]), .C(SLM_CLK_c), .D(n6909));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(pc_data_rx[2]), .C(SLM_CLK_c), .D(n6908));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(pc_data_rx[3]), .C(SLM_CLK_c), .D(n6907));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(pc_data_rx[4]), .C(SLM_CLK_c), .D(n6906));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(pc_data_rx[5]), .C(SLM_CLK_c), .D(n6905));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(pc_data_rx[6]), .C(SLM_CLK_c), .D(n6904));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(pc_data_rx[7]), .C(SLM_CLK_c), .D(n6903));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1607_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index_c[1]), 
            .I2(r_Bit_Index_c[2]), .I3(GND_net), .O(n340[2]));
    defparam i1607_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index_c[1]), 
            .I2(r_Bit_Index_c[2]), .I3(GND_net), .O(n9011));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_CARRY r_Clock_Count_1439_add_4_8 (.CI(n12192), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n12193));
    SB_LUT4 r_Clock_Count_1439_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n12191), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1439_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index_c[2]), .C(SLM_CLK_c), .E(n13008), 
            .D(n340[2]), .R(n13034));   // src/uart_rx.v(49[10] 144[8])
    SB_CARRY r_Clock_Count_1439_add_4_7 (.CI(n12191), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n12192));
    SB_LUT4 r_Clock_Count_1439_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n12190), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1439_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index_c[1]), .C(SLM_CLK_c), .E(n13008), 
            .D(n340[1]), .R(n13034));   // src/uart_rx.v(49[10] 144[8])
    SB_CARRY r_Clock_Count_1439_add_4_6 (.CI(n12190), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n12191));
    SB_LUT4 r_Clock_Count_1439_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n12189), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1439_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1439_add_4_5 (.CI(n12189), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n12190));
    SB_LUT4 r_Clock_Count_1439_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n12188), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1439_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1439_add_4_4 (.CI(n12188), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n12189));
    SB_LUT4 r_Clock_Count_1439_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n12187), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1439_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(SLM_CLK_c), .D(r_SM_Main_2__N_950[2]), 
            .R(n12875));   // src/uart_rx.v(49[10] 144[8])
    SB_CARRY r_Clock_Count_1439_add_4_3 (.CI(n12187), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n12188));
    SB_LUT4 r_Clock_Count_1439_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1439_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1439_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n12187));
    SB_DFFESR r_Clock_Count_1439__i9 (.Q(r_Clock_Count[9]), .C(SLM_CLK_c), 
            .E(n4913), .D(n45[9]), .R(n5532));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1439__i8 (.Q(r_Clock_Count[8]), .C(SLM_CLK_c), 
            .E(n4913), .D(n45[8]), .R(n5532));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1439__i7 (.Q(r_Clock_Count[7]), .C(SLM_CLK_c), 
            .E(n4913), .D(n45[7]), .R(n5532));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1439__i6 (.Q(r_Clock_Count[6]), .C(SLM_CLK_c), 
            .E(n4913), .D(n45[6]), .R(n5532));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1439__i5 (.Q(r_Clock_Count[5]), .C(SLM_CLK_c), 
            .E(n4913), .D(n45[5]), .R(n5532));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1439__i4 (.Q(r_Clock_Count[4]), .C(SLM_CLK_c), 
            .E(n4913), .D(n45[4]), .R(n5532));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1439__i0 (.Q(r_Clock_Count[0]), .C(SLM_CLK_c), 
            .E(n4913), .D(n45[0]), .R(n5532));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1439__i3 (.Q(r_Clock_Count[3]), .C(SLM_CLK_c), 
            .E(n4913), .D(n45[3]), .R(n5532));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1439__i2 (.Q(r_Clock_Count[2]), .C(SLM_CLK_c), 
            .E(n4913), .D(n45[2]), .R(n5532));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1439__i1 (.Q(r_Clock_Count[1]), .C(SLM_CLK_c), 
            .E(n4913), .D(n45[1]), .R(n5532));   // src/uart_rx.v(120[34:51])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(SLM_CLK_c), .D(n9053), 
            .R(r_SM_Main[2]));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(SLM_CLK_c), .D(UART_RX_c));   // src/uart_rx.v(41[10] 45[8])
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[4]), .I2(r_Clock_Count[3]), 
            .I3(n4691), .O(n8));   // src/uart_rx.v(68[17:52])
    defparam i3_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i4_3_lut (.I0(r_Clock_Count[1]), .I1(n8), .I2(r_Clock_Count[2]), 
            .I3(GND_net), .O(r_SM_Main_2__N_956[0]));   // src/uart_rx.v(68[17:52])
    defparam i4_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_77 (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[9]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_1399));   // src/uart_rx.v(68[17:52])
    defparam i1_2_lut_adj_77.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[7]), .I2(r_Clock_Count[5]), 
            .I3(n6_adj_1399), .O(n4691));   // src/uart_rx.v(68[17:52])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[1]), 
            .I3(GND_net), .O(n4_adj_1400));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7566_4_lut (.I0(r_Clock_Count[3]), .I1(n4691), .I2(r_Clock_Count[4]), 
            .I3(n4_adj_1400), .O(r_SM_Main_2__N_950[2]));
    defparam i7566_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n9011), .I1(r_SM_Main_2__N_950[2]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n9043));   // src/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_956[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // src/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i3_3_lut (.I0(n1), .I1(n9043), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // src/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index_c[2]), .I1(n4693), .I2(r_Bit_Index_c[1]), 
            .I3(GND_net), .O(n4787));
    defparam i2_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 equal_145_i4_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_9));   // src/uart_rx.v(97[17:39])
    defparam equal_145_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_148_i4_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_10));   // src/uart_rx.v(97[17:39])
    defparam equal_148_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_78 (.I0(n4693), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4794));   // src/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_78.LUT_INIT = 16'hbbbb;
    SB_LUT4 i12351_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n12875));   // src/uart_rx.v(52[7] 143[14])
    defparam i12351_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_950[2]), 
            .I3(r_SM_Main[0]), .O(n4870));   // src/uart_rx.v(52[7] 143[14])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n4870), 
            .I3(debug_led3), .O(n12411));   // src/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i12374_4_lut (.I0(r_SM_Main_2__N_950[2]), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n13008));
    defparam i12374_4_lut.LUT_INIT = 16'h0023;
    SB_LUT4 i12355_3_lut (.I0(n13008), .I1(n9011), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n13034));
    defparam i12355_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_950[2]), 
            .I2(r_SM_Main[1]), .I3(n4_adj_1398), .O(n9053));   // src/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h707a;
    SB_LUT4 i10915_2_lut_3_lut (.I0(r_SM_Main[0]), .I1(r_Rx_Data), .I2(r_SM_Main_2__N_956[0]), 
            .I3(GND_net), .O(n13024));
    defparam i10915_2_lut_3_lut.LUT_INIT = 16'ha8a8;
    
endmodule
//
// Verilog Description of module fifo_dc_32_lut_gen2
//

module fifo_dc_32_lut_gen2 (dc32_fifo_data_in, \REG.mem_1_9 , GND_net, 
            \REG.mem_6_9 , \REG.mem_7_9 , \REG.mem_4_9 , \REG.mem_5_9 , 
            \REG.mem_24_9 , \REG.mem_25_9 , \REG.mem_1_31 , \REG.mem_9_5 , 
            \REG.mem_8_5 , \REG.mem_26_9 , \REG.mem_27_9 , rd_grey_sync_r, 
            \REG.mem_17_25 , \REG.mem_6_16 , \REG.mem_7_16 , \REG.mem_1_7 , 
            \REG.mem_6_7 , \REG.mem_7_7 , \REG.mem_4_7 , \REG.mem_5_7 , 
            \REG.mem_10_23 , \REG.mem_11_23 , \REG.mem_5_16 , \REG.mem_4_16 , 
            \REG.mem_17_7 , \REG.mem_22_7 , \REG.mem_23_7 , \REG.mem_20_7 , 
            \REG.mem_21_7 , \REG.mem_9_23 , \REG.mem_8_23 , n7, n23, 
            FIFO_CLK_c, DEBUG_1_c, reset_per_frame, wr_fifo_en_w, \wr_addr_r[0] , 
            \REG.mem_22_29 , \REG.mem_23_29 , \REG.mem_21_29 , \REG.mem_20_29 , 
            DEBUG_5_c_0, SLM_CLK_c, \REG.mem_26_21 , \REG.mem_27_21 , 
            \REG.mem_26_25 , \REG.mem_27_25 , \REG.mem_25_25 , \REG.mem_24_25 , 
            \REG.mem_25_21 , \REG.mem_24_21 , \REG.mem_1_10 , \REG.mem_6_10 , 
            \REG.mem_7_10 , \REG.mem_4_10 , \REG.mem_5_10 , \REG.mem_1_26 , 
            n28, n12, dc32_fifo_empty, \wr_grey_sync_r[0] , \aempty_flag_impl.ae_flag_nxt_w , 
            dc32_fifo_almost_empty, n32, n16, \REG.mem_17_10 , \REG.mem_22_10 , 
            \REG.mem_23_10 , \REG.mem_20_10 , \REG.mem_21_10 , dc32_fifo_full, 
            \REG.mem_10_28 , \REG.mem_11_28 , \REG.mem_9_28 , \REG.mem_8_28 , 
            \REG.mem_17_29 , \rd_addr_nxt_c_5__N_573[3] , \rd_addr_nxt_c_5__N_573[1] , 
            n6, n22, \REG.mem_1_28 , \REG.mem_6_28 , \REG.mem_7_28 , 
            \REG.mem_4_28 , \REG.mem_5_28 , \REG.mem_1_2 , \REG.mem_6_2 , 
            \REG.mem_7_2 , \REG.mem_4_2 , \REG.mem_5_2 , \REG.mem_1_22 , 
            \REG.mem_6_22 , \REG.mem_7_22 , \REG.mem_4_22 , \REG.mem_5_22 , 
            \REG.mem_17_22 , \REG.mem_22_22 , \REG.mem_23_22 , \REG.mem_20_22 , 
            \REG.mem_21_22 , \rd_addr_nxt_c_5__N_573[4] , \REG.mem_5_18 , 
            \REG.mem_4_18 , \REG.mem_6_4 , \REG.mem_7_4 , \REG.mem_6_18 , 
            \REG.mem_7_18 , \REG.mem_10_8 , \REG.mem_11_8 , \REG.mem_9_8 , 
            \REG.mem_8_8 , \REG.mem_5_4 , \REG.mem_4_4 , \REG.mem_1_21 , 
            n7013, n7012, n7011, n7010, n7009, n7008, wp_sync1_r, 
            n7007, n7006, n7005, n7004, n7003, n7002, n7000, n6998, 
            n6997, n6996, n6995, n6994, n6993, rp_sync1_r, n6992, 
            n6991, n6990, n6989, \REG.mem_1_13 , n6930, n6928, \wr_addr_r[5] , 
            \REG.mem_6_30 , \REG.mem_7_30 , n6493, \REG.mem_27_31 , 
            n6492, \REG.mem_27_30 , n6491, \REG.mem_27_29 , n6490, 
            \REG.mem_27_28 , n6489, \REG.mem_27_27 , n6488, \REG.mem_27_26 , 
            n6487, n6486, \REG.mem_27_24 , n6485, \REG.mem_27_23 , 
            n6484, \REG.mem_27_22 , n6483, n6482, \REG.mem_27_20 , 
            n6481, \REG.mem_27_19 , n6480, \REG.mem_27_18 , n6479, 
            \REG.mem_27_17 , n6478, \REG.mem_27_16 , n6477, \REG.mem_27_15 , 
            n6476, \REG.mem_27_14 , n6475, \REG.mem_27_13 , n6474, 
            \REG.mem_27_12 , n6473, \REG.mem_27_11 , n6472, \REG.mem_27_10 , 
            n6471, n6470, \REG.mem_27_8 , n6469, \REG.mem_27_7 , n6468, 
            \REG.mem_27_6 , n6467, \REG.mem_27_5 , n6466, \REG.mem_27_4 , 
            n6465, \REG.mem_27_3 , n6464, \REG.mem_27_2 , n6463, \REG.mem_27_1 , 
            n6462, \REG.mem_27_0 , n6461, \REG.mem_26_31 , n6460, 
            \REG.mem_26_30 , n6459, \REG.mem_26_29 , n6458, \REG.mem_26_28 , 
            n6457, \REG.mem_26_27 , n6456, \REG.mem_26_26 , n6455, 
            n6454, \REG.mem_26_24 , n6453, \REG.mem_26_23 , n6452, 
            \REG.mem_26_22 , n6451, n6450, \REG.mem_26_20 , n6449, 
            \REG.mem_26_19 , n6448, \REG.mem_26_18 , n6447, \REG.mem_26_17 , 
            n6446, \REG.mem_26_16 , n6445, \REG.mem_26_15 , n6444, 
            \REG.mem_26_14 , n6443, \REG.mem_26_13 , n6442, \REG.mem_26_12 , 
            n6441, \REG.mem_26_11 , n6440, \REG.mem_26_10 , n6439, 
            n6438, \REG.mem_26_8 , n6437, \REG.mem_26_7 , n6436, \REG.mem_26_6 , 
            n6435, \REG.mem_26_5 , n6434, \REG.mem_26_4 , n6433, \REG.mem_26_3 , 
            n6432, \REG.mem_26_2 , n6431, \REG.mem_26_1 , n6430, \REG.mem_26_0 , 
            n6429, \REG.mem_25_31 , n6428, \REG.mem_25_30 , n6427, 
            \REG.mem_25_29 , n6426, \REG.mem_25_28 , n6425, \REG.mem_25_27 , 
            n6424, \REG.mem_25_26 , n6423, n6422, \REG.mem_25_24 , 
            n6421, \REG.mem_25_23 , n6420, \REG.mem_25_22 , n6419, 
            n6418, \REG.mem_25_20 , n6417, \REG.mem_25_19 , n6416, 
            \REG.mem_25_18 , n6415, \REG.mem_25_17 , n6414, \REG.mem_25_16 , 
            n6413, \REG.mem_25_15 , n6412, \REG.mem_25_14 , n6411, 
            \REG.mem_25_13 , n6410, \REG.mem_25_12 , n6409, \REG.mem_25_11 , 
            n6408, \REG.mem_25_10 , n6407, n6406, \REG.mem_25_8 , 
            n6405, \REG.mem_25_7 , n6404, \REG.mem_25_6 , n6403, \REG.mem_25_5 , 
            n6402, \REG.mem_25_4 , n6401, \REG.mem_25_3 , n6400, \REG.mem_25_2 , 
            n6399, \REG.mem_25_1 , n6398, \REG.mem_25_0 , n6397, \REG.mem_24_31 , 
            n6396, \REG.mem_24_30 , n6395, \REG.mem_24_29 , n6394, 
            \REG.mem_24_28 , n6393, \REG.mem_24_27 , n6392, \REG.mem_24_26 , 
            n6391, n6390, \REG.mem_24_24 , n6389, \REG.mem_24_23 , 
            n6388, \REG.mem_24_22 , n6387, n6386, \REG.mem_24_20 , 
            n6385, \REG.mem_24_19 , n6384, \REG.mem_24_18 , n6383, 
            \REG.mem_24_17 , n6382, \REG.mem_24_16 , n6381, \REG.mem_24_15 , 
            n6380, \REG.mem_24_14 , n6379, \REG.mem_24_13 , n6378, 
            \REG.mem_24_12 , n6377, \REG.mem_24_11 , n6376, \REG.mem_24_10 , 
            n6375, n6374, \REG.mem_24_8 , n6373, \REG.mem_24_7 , n6372, 
            \REG.mem_24_6 , n6371, \REG.mem_24_5 , n6370, \REG.mem_24_4 , 
            n6369, \REG.mem_24_3 , n6368, \REG.mem_24_2 , n6367, \REG.mem_24_1 , 
            n6366, \REG.mem_24_0 , n6365, \REG.mem_23_31 , n6364, 
            \REG.mem_23_30 , n6363, n6362, \REG.mem_23_28 , n6361, 
            \REG.mem_23_27 , n6360, \REG.mem_23_26 , n6359, \REG.mem_23_25 , 
            n6358, \REG.mem_23_24 , n6357, \REG.mem_23_23 , n6356, 
            n6355, \REG.mem_23_21 , n6354, \REG.mem_23_20 , n6353, 
            \REG.mem_23_19 , n6352, \REG.mem_23_18 , n6351, \REG.mem_23_17 , 
            n6350, \REG.mem_23_16 , n6349, \REG.mem_23_15 , n6348, 
            \REG.mem_23_14 , n6347, \REG.mem_23_13 , n6346, \REG.mem_23_12 , 
            n6345, \REG.mem_23_11 , n6344, n6343, \REG.mem_23_9 , 
            n6342, \REG.mem_23_8 , n6341, n6340, \REG.mem_23_6 , n6339, 
            \REG.mem_23_5 , n6338, \REG.mem_23_4 , n6337, \REG.mem_23_3 , 
            n6336, \REG.mem_23_2 , n6335, \REG.mem_23_1 , n6334, \REG.mem_23_0 , 
            n6333, \REG.mem_22_31 , n6332, \REG.mem_22_30 , n6331, 
            n6330, \REG.mem_22_28 , n6329, \REG.mem_22_27 , n6328, 
            \REG.mem_22_26 , n6327, \REG.mem_22_25 , n6326, \REG.mem_22_24 , 
            n6325, \REG.mem_22_23 , n6324, n6323, \REG.mem_22_21 , 
            n6322, \REG.mem_22_20 , n6321, \REG.mem_22_19 , n6320, 
            \REG.mem_22_18 , n6319, \REG.mem_22_17 , n6318, \REG.mem_22_16 , 
            n6317, \REG.mem_22_15 , n6316, \REG.mem_22_14 , n6315, 
            \REG.mem_22_13 , n6314, \REG.mem_22_12 , n6313, \REG.mem_22_11 , 
            n6312, n6311, \REG.mem_22_9 , n6310, \REG.mem_22_8 , n6309, 
            n6308, \REG.mem_22_6 , n6307, \REG.mem_22_5 , n6306, \REG.mem_22_4 , 
            n6305, \REG.mem_22_3 , n6304, \REG.mem_22_2 , n6303, \REG.mem_22_1 , 
            n6302, \REG.mem_22_0 , n6301, \REG.mem_21_31 , n6300, 
            \REG.mem_21_30 , n6299, n6298, \REG.mem_21_28 , n6297, 
            \REG.mem_21_27 , n6296, \REG.mem_21_26 , n6295, \REG.mem_21_25 , 
            n6294, \REG.mem_21_24 , n6293, \REG.mem_21_23 , n6292, 
            n6291, \REG.mem_21_21 , n6290, \REG.mem_21_20 , n6289, 
            \REG.mem_21_19 , n6288, \REG.mem_21_18 , n6287, \REG.mem_21_17 , 
            n6286, \REG.mem_21_16 , n6285, \REG.mem_21_15 , n6284, 
            \REG.mem_21_14 , n6283, \REG.mem_21_13 , n6282, \REG.mem_21_12 , 
            n6281, \REG.mem_21_11 , n6280, n6279, \REG.mem_21_9 , 
            n6278, \REG.mem_21_8 , n6277, n6276, \REG.mem_21_6 , n6275, 
            \REG.mem_21_5 , n6274, \REG.mem_21_4 , n6273, \REG.mem_21_3 , 
            n6272, \REG.mem_21_2 , n6271, \REG.mem_21_1 , n6270, \REG.mem_21_0 , 
            n6269, \REG.mem_20_31 , n6268, \REG.mem_20_30 , n6267, 
            n6266, \REG.mem_20_28 , n6265, \REG.mem_20_27 , n6264, 
            \REG.mem_20_26 , n6263, \REG.mem_20_25 , n6262, \REG.mem_20_24 , 
            n6261, \REG.mem_20_23 , n6260, n6259, \REG.mem_20_21 , 
            n6258, \REG.mem_20_20 , n6257, \REG.mem_20_19 , n6256, 
            \REG.mem_20_18 , n6255, \REG.mem_20_17 , n6254, \REG.mem_20_16 , 
            n6253, \REG.mem_20_15 , n6252, \REG.mem_20_14 , n6251, 
            \REG.mem_20_13 , n6250, \REG.mem_20_12 , n6249, \REG.mem_20_11 , 
            n6248, n6247, \REG.mem_20_9 , n6246, \REG.mem_20_8 , n6245, 
            n6244, \REG.mem_20_6 , n6243, \REG.mem_20_5 , n6242, \REG.mem_20_4 , 
            n6241, \REG.mem_20_3 , n6240, \REG.mem_20_2 , n6239, \REG.mem_20_1 , 
            n6238, \REG.mem_20_0 , n6173, \REG.mem_17_31 , n6172, 
            \REG.mem_17_30 , n6171, n6170, \REG.mem_17_28 , n6169, 
            \REG.mem_17_27 , n6168, \REG.mem_17_26 , n6167, n6166, 
            \REG.mem_17_24 , n6165, \REG.mem_17_23 , n6164, n6163, 
            \REG.mem_17_21 , n6162, \REG.mem_17_20 , n6161, \REG.mem_17_19 , 
            n6160, \REG.mem_17_18 , n6159, \REG.mem_17_17 , n6158, 
            \REG.mem_17_16 , n6157, \REG.mem_17_15 , n6156, \REG.mem_17_14 , 
            n6155, \REG.mem_17_13 , n6154, \REG.mem_17_12 , n6153, 
            \REG.mem_17_11 , n6152, n6151, \REG.mem_17_9 , n6150, 
            \REG.mem_17_8 , n6149, n6148, \REG.mem_17_6 , n6147, \REG.mem_17_5 , 
            n6146, \REG.mem_17_4 , n6145, \REG.mem_17_3 , n6144, \REG.mem_17_2 , 
            n6143, \REG.mem_17_1 , n6142, \REG.mem_17_0 , \REG.mem_5_30 , 
            \REG.mem_4_30 , \REG.mem_1_1 , \REG.mem_6_1 , \REG.mem_7_1 , 
            \REG.mem_4_1 , \REG.mem_5_1 , \REG.mem_6_21 , \REG.mem_7_21 , 
            \REG.mem_5_21 , \REG.mem_4_21 , \REG.mem_1_30 , \REG.mem_10_21 , 
            \REG.mem_11_21 , \REG.mem_1_19 , \REG.mem_6_19 , \REG.mem_7_19 , 
            \REG.mem_5_19 , \REG.mem_4_19 , \REG.mem_9_21 , \REG.mem_8_21 , 
            \wr_addr_p1_w[0] , \REG.mem_6_13 , \REG.mem_7_13 , \REG.mem_5_13 , 
            \REG.mem_4_13 , \REG.mem_10_13 , \REG.mem_11_13 , \REG.mem_9_13 , 
            \REG.mem_8_13 , \REG.mem_10_19 , \REG.mem_11_19 , \REG.mem_9_19 , 
            \REG.mem_8_19 , \REG.mem_1_27 , \REG.mem_6_27 , \REG.mem_7_27 , 
            \REG.mem_4_27 , \REG.mem_5_27 , \REG.mem_1_6 , \REG.mem_8_2 , 
            \REG.mem_9_2 , \REG.mem_10_2 , \REG.mem_11_2 , \wr_addr_nxt_c[2] , 
            VCC_net, dc32_fifo_write_enable, \REG.mem_1_0 , \REG.mem_10_15 , 
            \REG.mem_11_15 , \REG.mem_9_15 , \REG.mem_8_15 , \dc32_fifo_data_out[1] , 
            \REG.mem_10_11 , \REG.mem_11_11 , \REG.mem_9_11 , \REG.mem_8_11 , 
            \dc32_fifo_data_out[2] , \dc32_fifo_data_out[3] , \dc32_fifo_data_out[4] , 
            \dc32_fifo_data_out[5] , \dc32_fifo_data_out[6] , \dc32_fifo_data_out[7] , 
            \dc32_fifo_data_out[8] , \dc32_fifo_data_out[9] , \dc32_fifo_data_out[10] , 
            \dc32_fifo_data_out[11] , \dc32_fifo_data_out[12] , \dc32_fifo_data_out[13] , 
            \dc32_fifo_data_out[14] , \dc32_fifo_data_out[15] , \dc32_fifo_data_out[16] , 
            \dc32_fifo_data_out[17] , \dc32_fifo_data_out[18] , \dc32_fifo_data_out[19] , 
            \dc32_fifo_data_out[20] , \dc32_fifo_data_out[21] , \dc32_fifo_data_out[22] , 
            \dc32_fifo_data_out[23] , \dc32_fifo_data_out[24] , \dc32_fifo_data_out[25] , 
            \dc32_fifo_data_out[26] , \dc32_fifo_data_out[27] , \dc32_fifo_data_out[28] , 
            \dc32_fifo_data_out[29] , \dc32_fifo_data_out[30] , \dc32_fifo_data_out[31] , 
            n7_adj_6, n8, n25, n5981, \REG.mem_11_31 , \REG.mem_1_23 , 
            n5980, \REG.mem_11_30 , \REG.mem_6_6 , \REG.mem_7_6 , \REG.mem_5_6 , 
            \REG.mem_4_6 , n5979, \REG.mem_11_29 , \REG.mem_10_29 , 
            n5978, n5977, \REG.mem_11_27 , n5976, \REG.mem_11_26 , 
            n5975, \REG.mem_11_25 , n5974, \REG.mem_11_24 , \REG.mem_9_29 , 
            \REG.mem_8_29 , n5973, n5972, \REG.mem_11_22 , n29, \REG.mem_8_17 , 
            \REG.mem_9_17 , \REG.mem_10_17 , \REG.mem_11_17 , \REG.mem_1_24 , 
            n5971, n5970, \REG.mem_11_20 , \REG.mem_6_31 , \REG.mem_7_31 , 
            \REG.mem_5_31 , \REG.mem_4_31 , \wr_grey_sync_r[1] , n24, 
            n13, n8_adj_7, \REG.mem_6_23 , \REG.mem_7_23 , \REG.mem_5_23 , 
            \REG.mem_4_23 , \REG.mem_10_6 , \REG.mem_11_6 , n5969, \REG.mem_9_6 , 
            \REG.mem_8_6 , \wr_grey_sync_r[2] , \wr_grey_sync_r[3] , \wr_grey_sync_r[4] , 
            n5968, \REG.mem_11_18 , n5967, n5966, \REG.mem_11_16 , 
            n5965, n5964, \REG.mem_11_14 , n5963, n5962, \REG.mem_11_12 , 
            n5961, n5960, \REG.mem_11_10 , n5959, \REG.mem_11_9 , 
            n5958, n5957, \REG.mem_11_7 , n5956, n5955, \REG.mem_11_5 , 
            n5954, \REG.mem_11_4 , n5953, \REG.mem_11_3 , \REG.mem_10_22 , 
            n5952, n5951, \REG.mem_11_1 , n5950, \REG.mem_11_0 , n5949, 
            \REG.mem_10_31 , n5948, \REG.mem_10_30 , n5947, n5946, 
            n5945, \REG.mem_10_27 , \REG.mem_9_22 , \REG.mem_8_22 , 
            n5944, \REG.mem_10_26 , \REG.mem_1_18 , n5943, \REG.mem_10_25 , 
            n5942, \REG.mem_10_24 , n5611, \REG.mem_6_24 , \REG.mem_7_24 , 
            \REG.mem_5_24 , \REG.mem_4_24 , \REG.mem_1_4 , \REG.mem_9_24 , 
            \REG.mem_8_24 , \REG.mem_6_0 , \REG.mem_7_0 , \REG.mem_5_0 , 
            \REG.mem_4_0 , \REG.mem_10_4 , n5610, n5941, n5940, n5939, 
            n5938, \REG.mem_10_20 , n5937, n5608, n5604, n5603, 
            n5602, n5936, \REG.mem_10_18 , n5935, n5934, \REG.mem_10_16 , 
            n5933, \REG.mem_1_17 , \REG.mem_9_4 , \REG.mem_8_4 , \REG.mem_6_17 , 
            \REG.mem_7_17 , \REG.mem_4_17 , \REG.mem_5_17 , dc32_fifo_read_enable, 
            n5932, \REG.mem_10_14 , n5931, n5930, \REG.mem_10_12 , 
            n5929, n5928, \REG.mem_10_10 , n5927, \REG.mem_10_9 , 
            n5926, n5925, \REG.mem_10_7 , n5924, n5923, \REG.mem_10_5 , 
            n5922, n5921, \REG.mem_10_3 , n5920, n5919, \REG.mem_10_1 , 
            n5918, \REG.mem_10_0 , n5917, \REG.mem_9_31 , n5916, \REG.mem_9_30 , 
            n5915, n5914, n5913, \REG.mem_9_27 , n5912, \REG.mem_9_26 , 
            n5911, \REG.mem_9_25 , n5910, n5909, n5908, n5907, n5906, 
            \REG.mem_9_20 , n5905, n5904, \REG.mem_9_18 , n5903, n5902, 
            \REG.mem_9_16 , n5901, n5900, \REG.mem_9_14 , n5899, n5898, 
            \REG.mem_9_12 , n5897, n5896, \REG.mem_9_10 , n5895, \REG.mem_9_9 , 
            n5894, n5893, \REG.mem_9_7 , n5892, n5891, n5890, n5889, 
            \REG.mem_9_3 , n5888, n5887, \REG.mem_9_1 , n5886, \REG.mem_9_0 , 
            n5885, \REG.mem_8_31 , n5884, \REG.mem_8_30 , n5883, n5882, 
            n5881, \REG.mem_8_27 , n5880, \REG.mem_8_26 , n5879, \REG.mem_8_25 , 
            n5878, n5877, n5876, n5875, n5874, \REG.mem_8_20 , n5873, 
            n5872, \REG.mem_8_18 , n5871, n5870, \REG.mem_8_16 , n5869, 
            n5868, \REG.mem_8_14 , n5867, n5866, \REG.mem_8_12 , n5865, 
            n5864, \REG.mem_8_10 , n5863, \REG.mem_8_9 , n5862, n5861, 
            \REG.mem_8_7 , n5860, n5859, n5858, n5857, \REG.mem_8_3 , 
            n5856, n5855, \REG.mem_8_1 , n5854, \REG.mem_8_0 , n5853, 
            n5852, n5851, \REG.mem_7_29 , n5850, n5849, n5848, \REG.mem_7_26 , 
            n5847, \REG.mem_7_25 , n5846, n5845, n5844, n5843, n5842, 
            \REG.mem_7_20 , n5841, n5840, n5839, n5838, n5837, \REG.mem_7_15 , 
            n5836, \REG.mem_7_14 , n5835, n5834, \REG.mem_7_12 , n5833, 
            \REG.mem_7_11 , n5832, n5831, n5830, \REG.mem_7_8 , n5829, 
            n5828, n5827, \REG.mem_7_5 , n5826, n5825, \REG.mem_7_3 , 
            n5824, n5823, n5822, n5821, n5820, n5819, \REG.mem_6_29 , 
            n5818, n5817, n5816, \REG.mem_6_26 , n5815, \REG.mem_6_25 , 
            n5814, n5813, n5812, n5811, n5810, \REG.mem_6_20 , n5809, 
            n5808, n5807, n5806, n5805, \REG.mem_6_15 , n5804, \REG.mem_6_14 , 
            n5803, n5802, \REG.mem_6_12 , n5801, \REG.mem_6_11 , n5800, 
            n5799, n5798, \REG.mem_6_8 , n5797, n5796, n5795, \REG.mem_6_5 , 
            n5794, n5793, \REG.mem_6_3 , n5792, n5791, n5790, n5789, 
            n5788, n5600, \REG.mem_1_3 , n5787, \REG.mem_5_29 , n25_adj_8, 
            n9, n5786, n5785, n5784, \REG.mem_5_26 , n5783, \REG.mem_5_25 , 
            n5782, \REG.mem_1_16 , n5781, n5780, n5779, n5778, \REG.mem_5_20 , 
            n5777, n5776, n5775, n5774, n5773, \REG.mem_5_15 , n5772, 
            \REG.mem_5_14 , n5771, n5770, \REG.mem_5_12 , n5769, \REG.mem_5_11 , 
            \REG.mem_1_25 , n5768, n5767, n5766, \REG.mem_5_8 , n5765, 
            n10, n26, n5596, n5764, n5595, \REG.mem_1_5 , n5594, 
            n5593, n5590, n5589, n5588, n5587, n5763, \REG.mem_5_5 , 
            \REG.mem_4_26 , n5762, n5761, \REG.mem_5_3 , n5760, n5759, 
            n5586, n5758, n5757, n5756, n5755, \REG.mem_4_29 , \wr_addr_nxt_c[4] , 
            n5754, n5753, n5752, n5751, \REG.mem_4_25 , n5750, n5749, 
            n5748, n5747, n5585, \REG.mem_1_29 , n5583, n5582, n5581, 
            \REG.mem_1_8 , n5580, n5577, n5746, \REG.mem_4_20 , n5745, 
            n5744, n5743, n5742, n5741, \REG.mem_4_15 , n5740, \REG.mem_4_14 , 
            n5739, n5738, \REG.mem_4_12 , n5574, n5572, n5571, \REG.mem_1_11 , 
            n5737, \REG.mem_4_11 , n5736, n5735, n5734, \REG.mem_4_8 , 
            n5733, n5732, n5731, \REG.mem_4_5 , n5730, n5729, \REG.mem_4_3 , 
            n5567, n5565, \REG.mem_1_20 , n5564, \REG.mem_1_12 , n5560, 
            n5559, \REG.mem_1_14 , n5558, \REG.mem_1_15 , n5557, n5556, 
            n5555, n5554, n5551, n5550, n5728, n5727, n5726, n11, 
            n27) /* synthesis syn_module_defined=1 */ ;
    input [31:0]dc32_fifo_data_in;
    output \REG.mem_1_9 ;
    input GND_net;
    output \REG.mem_6_9 ;
    output \REG.mem_7_9 ;
    output \REG.mem_4_9 ;
    output \REG.mem_5_9 ;
    output \REG.mem_24_9 ;
    output \REG.mem_25_9 ;
    output \REG.mem_1_31 ;
    output \REG.mem_9_5 ;
    output \REG.mem_8_5 ;
    output \REG.mem_26_9 ;
    output \REG.mem_27_9 ;
    output [5:0]rd_grey_sync_r;
    output \REG.mem_17_25 ;
    output \REG.mem_6_16 ;
    output \REG.mem_7_16 ;
    output \REG.mem_1_7 ;
    output \REG.mem_6_7 ;
    output \REG.mem_7_7 ;
    output \REG.mem_4_7 ;
    output \REG.mem_5_7 ;
    output \REG.mem_10_23 ;
    output \REG.mem_11_23 ;
    output \REG.mem_5_16 ;
    output \REG.mem_4_16 ;
    output \REG.mem_17_7 ;
    output \REG.mem_22_7 ;
    output \REG.mem_23_7 ;
    output \REG.mem_20_7 ;
    output \REG.mem_21_7 ;
    output \REG.mem_9_23 ;
    output \REG.mem_8_23 ;
    output n7;
    output n23;
    input FIFO_CLK_c;
    output DEBUG_1_c;
    input reset_per_frame;
    output wr_fifo_en_w;
    output \wr_addr_r[0] ;
    output \REG.mem_22_29 ;
    output \REG.mem_23_29 ;
    output \REG.mem_21_29 ;
    output \REG.mem_20_29 ;
    output DEBUG_5_c_0;
    input SLM_CLK_c;
    output \REG.mem_26_21 ;
    output \REG.mem_27_21 ;
    output \REG.mem_26_25 ;
    output \REG.mem_27_25 ;
    output \REG.mem_25_25 ;
    output \REG.mem_24_25 ;
    output \REG.mem_25_21 ;
    output \REG.mem_24_21 ;
    output \REG.mem_1_10 ;
    output \REG.mem_6_10 ;
    output \REG.mem_7_10 ;
    output \REG.mem_4_10 ;
    output \REG.mem_5_10 ;
    output \REG.mem_1_26 ;
    output n28;
    output n12;
    output dc32_fifo_empty;
    output \wr_grey_sync_r[0] ;
    input \aempty_flag_impl.ae_flag_nxt_w ;
    output dc32_fifo_almost_empty;
    output n32;
    output n16;
    output \REG.mem_17_10 ;
    output \REG.mem_22_10 ;
    output \REG.mem_23_10 ;
    output \REG.mem_20_10 ;
    output \REG.mem_21_10 ;
    output dc32_fifo_full;
    output \REG.mem_10_28 ;
    output \REG.mem_11_28 ;
    output \REG.mem_9_28 ;
    output \REG.mem_8_28 ;
    output \REG.mem_17_29 ;
    output \rd_addr_nxt_c_5__N_573[3] ;
    output \rd_addr_nxt_c_5__N_573[1] ;
    output n6;
    output n22;
    output \REG.mem_1_28 ;
    output \REG.mem_6_28 ;
    output \REG.mem_7_28 ;
    output \REG.mem_4_28 ;
    output \REG.mem_5_28 ;
    output \REG.mem_1_2 ;
    output \REG.mem_6_2 ;
    output \REG.mem_7_2 ;
    output \REG.mem_4_2 ;
    output \REG.mem_5_2 ;
    output \REG.mem_1_22 ;
    output \REG.mem_6_22 ;
    output \REG.mem_7_22 ;
    output \REG.mem_4_22 ;
    output \REG.mem_5_22 ;
    output \REG.mem_17_22 ;
    output \REG.mem_22_22 ;
    output \REG.mem_23_22 ;
    output \REG.mem_20_22 ;
    output \REG.mem_21_22 ;
    output \rd_addr_nxt_c_5__N_573[4] ;
    output \REG.mem_5_18 ;
    output \REG.mem_4_18 ;
    output \REG.mem_6_4 ;
    output \REG.mem_7_4 ;
    output \REG.mem_6_18 ;
    output \REG.mem_7_18 ;
    output \REG.mem_10_8 ;
    output \REG.mem_11_8 ;
    output \REG.mem_9_8 ;
    output \REG.mem_8_8 ;
    output \REG.mem_5_4 ;
    output \REG.mem_4_4 ;
    output \REG.mem_1_21 ;
    input n7013;
    input n7012;
    input n7011;
    input n7010;
    input n7009;
    input n7008;
    output [5:0]wp_sync1_r;
    input n7007;
    input n7006;
    input n7005;
    input n7004;
    input n7003;
    input n7002;
    input n7000;
    input n6998;
    input n6997;
    input n6996;
    input n6995;
    input n6994;
    input n6993;
    output [5:0]rp_sync1_r;
    input n6992;
    input n6991;
    input n6990;
    input n6989;
    output \REG.mem_1_13 ;
    input n6930;
    input n6928;
    output \wr_addr_r[5] ;
    output \REG.mem_6_30 ;
    output \REG.mem_7_30 ;
    input n6493;
    output \REG.mem_27_31 ;
    input n6492;
    output \REG.mem_27_30 ;
    input n6491;
    output \REG.mem_27_29 ;
    input n6490;
    output \REG.mem_27_28 ;
    input n6489;
    output \REG.mem_27_27 ;
    input n6488;
    output \REG.mem_27_26 ;
    input n6487;
    input n6486;
    output \REG.mem_27_24 ;
    input n6485;
    output \REG.mem_27_23 ;
    input n6484;
    output \REG.mem_27_22 ;
    input n6483;
    input n6482;
    output \REG.mem_27_20 ;
    input n6481;
    output \REG.mem_27_19 ;
    input n6480;
    output \REG.mem_27_18 ;
    input n6479;
    output \REG.mem_27_17 ;
    input n6478;
    output \REG.mem_27_16 ;
    input n6477;
    output \REG.mem_27_15 ;
    input n6476;
    output \REG.mem_27_14 ;
    input n6475;
    output \REG.mem_27_13 ;
    input n6474;
    output \REG.mem_27_12 ;
    input n6473;
    output \REG.mem_27_11 ;
    input n6472;
    output \REG.mem_27_10 ;
    input n6471;
    input n6470;
    output \REG.mem_27_8 ;
    input n6469;
    output \REG.mem_27_7 ;
    input n6468;
    output \REG.mem_27_6 ;
    input n6467;
    output \REG.mem_27_5 ;
    input n6466;
    output \REG.mem_27_4 ;
    input n6465;
    output \REG.mem_27_3 ;
    input n6464;
    output \REG.mem_27_2 ;
    input n6463;
    output \REG.mem_27_1 ;
    input n6462;
    output \REG.mem_27_0 ;
    input n6461;
    output \REG.mem_26_31 ;
    input n6460;
    output \REG.mem_26_30 ;
    input n6459;
    output \REG.mem_26_29 ;
    input n6458;
    output \REG.mem_26_28 ;
    input n6457;
    output \REG.mem_26_27 ;
    input n6456;
    output \REG.mem_26_26 ;
    input n6455;
    input n6454;
    output \REG.mem_26_24 ;
    input n6453;
    output \REG.mem_26_23 ;
    input n6452;
    output \REG.mem_26_22 ;
    input n6451;
    input n6450;
    output \REG.mem_26_20 ;
    input n6449;
    output \REG.mem_26_19 ;
    input n6448;
    output \REG.mem_26_18 ;
    input n6447;
    output \REG.mem_26_17 ;
    input n6446;
    output \REG.mem_26_16 ;
    input n6445;
    output \REG.mem_26_15 ;
    input n6444;
    output \REG.mem_26_14 ;
    input n6443;
    output \REG.mem_26_13 ;
    input n6442;
    output \REG.mem_26_12 ;
    input n6441;
    output \REG.mem_26_11 ;
    input n6440;
    output \REG.mem_26_10 ;
    input n6439;
    input n6438;
    output \REG.mem_26_8 ;
    input n6437;
    output \REG.mem_26_7 ;
    input n6436;
    output \REG.mem_26_6 ;
    input n6435;
    output \REG.mem_26_5 ;
    input n6434;
    output \REG.mem_26_4 ;
    input n6433;
    output \REG.mem_26_3 ;
    input n6432;
    output \REG.mem_26_2 ;
    input n6431;
    output \REG.mem_26_1 ;
    input n6430;
    output \REG.mem_26_0 ;
    input n6429;
    output \REG.mem_25_31 ;
    input n6428;
    output \REG.mem_25_30 ;
    input n6427;
    output \REG.mem_25_29 ;
    input n6426;
    output \REG.mem_25_28 ;
    input n6425;
    output \REG.mem_25_27 ;
    input n6424;
    output \REG.mem_25_26 ;
    input n6423;
    input n6422;
    output \REG.mem_25_24 ;
    input n6421;
    output \REG.mem_25_23 ;
    input n6420;
    output \REG.mem_25_22 ;
    input n6419;
    input n6418;
    output \REG.mem_25_20 ;
    input n6417;
    output \REG.mem_25_19 ;
    input n6416;
    output \REG.mem_25_18 ;
    input n6415;
    output \REG.mem_25_17 ;
    input n6414;
    output \REG.mem_25_16 ;
    input n6413;
    output \REG.mem_25_15 ;
    input n6412;
    output \REG.mem_25_14 ;
    input n6411;
    output \REG.mem_25_13 ;
    input n6410;
    output \REG.mem_25_12 ;
    input n6409;
    output \REG.mem_25_11 ;
    input n6408;
    output \REG.mem_25_10 ;
    input n6407;
    input n6406;
    output \REG.mem_25_8 ;
    input n6405;
    output \REG.mem_25_7 ;
    input n6404;
    output \REG.mem_25_6 ;
    input n6403;
    output \REG.mem_25_5 ;
    input n6402;
    output \REG.mem_25_4 ;
    input n6401;
    output \REG.mem_25_3 ;
    input n6400;
    output \REG.mem_25_2 ;
    input n6399;
    output \REG.mem_25_1 ;
    input n6398;
    output \REG.mem_25_0 ;
    input n6397;
    output \REG.mem_24_31 ;
    input n6396;
    output \REG.mem_24_30 ;
    input n6395;
    output \REG.mem_24_29 ;
    input n6394;
    output \REG.mem_24_28 ;
    input n6393;
    output \REG.mem_24_27 ;
    input n6392;
    output \REG.mem_24_26 ;
    input n6391;
    input n6390;
    output \REG.mem_24_24 ;
    input n6389;
    output \REG.mem_24_23 ;
    input n6388;
    output \REG.mem_24_22 ;
    input n6387;
    input n6386;
    output \REG.mem_24_20 ;
    input n6385;
    output \REG.mem_24_19 ;
    input n6384;
    output \REG.mem_24_18 ;
    input n6383;
    output \REG.mem_24_17 ;
    input n6382;
    output \REG.mem_24_16 ;
    input n6381;
    output \REG.mem_24_15 ;
    input n6380;
    output \REG.mem_24_14 ;
    input n6379;
    output \REG.mem_24_13 ;
    input n6378;
    output \REG.mem_24_12 ;
    input n6377;
    output \REG.mem_24_11 ;
    input n6376;
    output \REG.mem_24_10 ;
    input n6375;
    input n6374;
    output \REG.mem_24_8 ;
    input n6373;
    output \REG.mem_24_7 ;
    input n6372;
    output \REG.mem_24_6 ;
    input n6371;
    output \REG.mem_24_5 ;
    input n6370;
    output \REG.mem_24_4 ;
    input n6369;
    output \REG.mem_24_3 ;
    input n6368;
    output \REG.mem_24_2 ;
    input n6367;
    output \REG.mem_24_1 ;
    input n6366;
    output \REG.mem_24_0 ;
    input n6365;
    output \REG.mem_23_31 ;
    input n6364;
    output \REG.mem_23_30 ;
    input n6363;
    input n6362;
    output \REG.mem_23_28 ;
    input n6361;
    output \REG.mem_23_27 ;
    input n6360;
    output \REG.mem_23_26 ;
    input n6359;
    output \REG.mem_23_25 ;
    input n6358;
    output \REG.mem_23_24 ;
    input n6357;
    output \REG.mem_23_23 ;
    input n6356;
    input n6355;
    output \REG.mem_23_21 ;
    input n6354;
    output \REG.mem_23_20 ;
    input n6353;
    output \REG.mem_23_19 ;
    input n6352;
    output \REG.mem_23_18 ;
    input n6351;
    output \REG.mem_23_17 ;
    input n6350;
    output \REG.mem_23_16 ;
    input n6349;
    output \REG.mem_23_15 ;
    input n6348;
    output \REG.mem_23_14 ;
    input n6347;
    output \REG.mem_23_13 ;
    input n6346;
    output \REG.mem_23_12 ;
    input n6345;
    output \REG.mem_23_11 ;
    input n6344;
    input n6343;
    output \REG.mem_23_9 ;
    input n6342;
    output \REG.mem_23_8 ;
    input n6341;
    input n6340;
    output \REG.mem_23_6 ;
    input n6339;
    output \REG.mem_23_5 ;
    input n6338;
    output \REG.mem_23_4 ;
    input n6337;
    output \REG.mem_23_3 ;
    input n6336;
    output \REG.mem_23_2 ;
    input n6335;
    output \REG.mem_23_1 ;
    input n6334;
    output \REG.mem_23_0 ;
    input n6333;
    output \REG.mem_22_31 ;
    input n6332;
    output \REG.mem_22_30 ;
    input n6331;
    input n6330;
    output \REG.mem_22_28 ;
    input n6329;
    output \REG.mem_22_27 ;
    input n6328;
    output \REG.mem_22_26 ;
    input n6327;
    output \REG.mem_22_25 ;
    input n6326;
    output \REG.mem_22_24 ;
    input n6325;
    output \REG.mem_22_23 ;
    input n6324;
    input n6323;
    output \REG.mem_22_21 ;
    input n6322;
    output \REG.mem_22_20 ;
    input n6321;
    output \REG.mem_22_19 ;
    input n6320;
    output \REG.mem_22_18 ;
    input n6319;
    output \REG.mem_22_17 ;
    input n6318;
    output \REG.mem_22_16 ;
    input n6317;
    output \REG.mem_22_15 ;
    input n6316;
    output \REG.mem_22_14 ;
    input n6315;
    output \REG.mem_22_13 ;
    input n6314;
    output \REG.mem_22_12 ;
    input n6313;
    output \REG.mem_22_11 ;
    input n6312;
    input n6311;
    output \REG.mem_22_9 ;
    input n6310;
    output \REG.mem_22_8 ;
    input n6309;
    input n6308;
    output \REG.mem_22_6 ;
    input n6307;
    output \REG.mem_22_5 ;
    input n6306;
    output \REG.mem_22_4 ;
    input n6305;
    output \REG.mem_22_3 ;
    input n6304;
    output \REG.mem_22_2 ;
    input n6303;
    output \REG.mem_22_1 ;
    input n6302;
    output \REG.mem_22_0 ;
    input n6301;
    output \REG.mem_21_31 ;
    input n6300;
    output \REG.mem_21_30 ;
    input n6299;
    input n6298;
    output \REG.mem_21_28 ;
    input n6297;
    output \REG.mem_21_27 ;
    input n6296;
    output \REG.mem_21_26 ;
    input n6295;
    output \REG.mem_21_25 ;
    input n6294;
    output \REG.mem_21_24 ;
    input n6293;
    output \REG.mem_21_23 ;
    input n6292;
    input n6291;
    output \REG.mem_21_21 ;
    input n6290;
    output \REG.mem_21_20 ;
    input n6289;
    output \REG.mem_21_19 ;
    input n6288;
    output \REG.mem_21_18 ;
    input n6287;
    output \REG.mem_21_17 ;
    input n6286;
    output \REG.mem_21_16 ;
    input n6285;
    output \REG.mem_21_15 ;
    input n6284;
    output \REG.mem_21_14 ;
    input n6283;
    output \REG.mem_21_13 ;
    input n6282;
    output \REG.mem_21_12 ;
    input n6281;
    output \REG.mem_21_11 ;
    input n6280;
    input n6279;
    output \REG.mem_21_9 ;
    input n6278;
    output \REG.mem_21_8 ;
    input n6277;
    input n6276;
    output \REG.mem_21_6 ;
    input n6275;
    output \REG.mem_21_5 ;
    input n6274;
    output \REG.mem_21_4 ;
    input n6273;
    output \REG.mem_21_3 ;
    input n6272;
    output \REG.mem_21_2 ;
    input n6271;
    output \REG.mem_21_1 ;
    input n6270;
    output \REG.mem_21_0 ;
    input n6269;
    output \REG.mem_20_31 ;
    input n6268;
    output \REG.mem_20_30 ;
    input n6267;
    input n6266;
    output \REG.mem_20_28 ;
    input n6265;
    output \REG.mem_20_27 ;
    input n6264;
    output \REG.mem_20_26 ;
    input n6263;
    output \REG.mem_20_25 ;
    input n6262;
    output \REG.mem_20_24 ;
    input n6261;
    output \REG.mem_20_23 ;
    input n6260;
    input n6259;
    output \REG.mem_20_21 ;
    input n6258;
    output \REG.mem_20_20 ;
    input n6257;
    output \REG.mem_20_19 ;
    input n6256;
    output \REG.mem_20_18 ;
    input n6255;
    output \REG.mem_20_17 ;
    input n6254;
    output \REG.mem_20_16 ;
    input n6253;
    output \REG.mem_20_15 ;
    input n6252;
    output \REG.mem_20_14 ;
    input n6251;
    output \REG.mem_20_13 ;
    input n6250;
    output \REG.mem_20_12 ;
    input n6249;
    output \REG.mem_20_11 ;
    input n6248;
    input n6247;
    output \REG.mem_20_9 ;
    input n6246;
    output \REG.mem_20_8 ;
    input n6245;
    input n6244;
    output \REG.mem_20_6 ;
    input n6243;
    output \REG.mem_20_5 ;
    input n6242;
    output \REG.mem_20_4 ;
    input n6241;
    output \REG.mem_20_3 ;
    input n6240;
    output \REG.mem_20_2 ;
    input n6239;
    output \REG.mem_20_1 ;
    input n6238;
    output \REG.mem_20_0 ;
    input n6173;
    output \REG.mem_17_31 ;
    input n6172;
    output \REG.mem_17_30 ;
    input n6171;
    input n6170;
    output \REG.mem_17_28 ;
    input n6169;
    output \REG.mem_17_27 ;
    input n6168;
    output \REG.mem_17_26 ;
    input n6167;
    input n6166;
    output \REG.mem_17_24 ;
    input n6165;
    output \REG.mem_17_23 ;
    input n6164;
    input n6163;
    output \REG.mem_17_21 ;
    input n6162;
    output \REG.mem_17_20 ;
    input n6161;
    output \REG.mem_17_19 ;
    input n6160;
    output \REG.mem_17_18 ;
    input n6159;
    output \REG.mem_17_17 ;
    input n6158;
    output \REG.mem_17_16 ;
    input n6157;
    output \REG.mem_17_15 ;
    input n6156;
    output \REG.mem_17_14 ;
    input n6155;
    output \REG.mem_17_13 ;
    input n6154;
    output \REG.mem_17_12 ;
    input n6153;
    output \REG.mem_17_11 ;
    input n6152;
    input n6151;
    output \REG.mem_17_9 ;
    input n6150;
    output \REG.mem_17_8 ;
    input n6149;
    input n6148;
    output \REG.mem_17_6 ;
    input n6147;
    output \REG.mem_17_5 ;
    input n6146;
    output \REG.mem_17_4 ;
    input n6145;
    output \REG.mem_17_3 ;
    input n6144;
    output \REG.mem_17_2 ;
    input n6143;
    output \REG.mem_17_1 ;
    input n6142;
    output \REG.mem_17_0 ;
    output \REG.mem_5_30 ;
    output \REG.mem_4_30 ;
    output \REG.mem_1_1 ;
    output \REG.mem_6_1 ;
    output \REG.mem_7_1 ;
    output \REG.mem_4_1 ;
    output \REG.mem_5_1 ;
    output \REG.mem_6_21 ;
    output \REG.mem_7_21 ;
    output \REG.mem_5_21 ;
    output \REG.mem_4_21 ;
    output \REG.mem_1_30 ;
    output \REG.mem_10_21 ;
    output \REG.mem_11_21 ;
    output \REG.mem_1_19 ;
    output \REG.mem_6_19 ;
    output \REG.mem_7_19 ;
    output \REG.mem_5_19 ;
    output \REG.mem_4_19 ;
    output \REG.mem_9_21 ;
    output \REG.mem_8_21 ;
    output \wr_addr_p1_w[0] ;
    output \REG.mem_6_13 ;
    output \REG.mem_7_13 ;
    output \REG.mem_5_13 ;
    output \REG.mem_4_13 ;
    output \REG.mem_10_13 ;
    output \REG.mem_11_13 ;
    output \REG.mem_9_13 ;
    output \REG.mem_8_13 ;
    output \REG.mem_10_19 ;
    output \REG.mem_11_19 ;
    output \REG.mem_9_19 ;
    output \REG.mem_8_19 ;
    output \REG.mem_1_27 ;
    output \REG.mem_6_27 ;
    output \REG.mem_7_27 ;
    output \REG.mem_4_27 ;
    output \REG.mem_5_27 ;
    output \REG.mem_1_6 ;
    output \REG.mem_8_2 ;
    output \REG.mem_9_2 ;
    output \REG.mem_10_2 ;
    output \REG.mem_11_2 ;
    output \wr_addr_nxt_c[2] ;
    input VCC_net;
    input dc32_fifo_write_enable;
    output \REG.mem_1_0 ;
    output \REG.mem_10_15 ;
    output \REG.mem_11_15 ;
    output \REG.mem_9_15 ;
    output \REG.mem_8_15 ;
    output \dc32_fifo_data_out[1] ;
    output \REG.mem_10_11 ;
    output \REG.mem_11_11 ;
    output \REG.mem_9_11 ;
    output \REG.mem_8_11 ;
    output \dc32_fifo_data_out[2] ;
    output \dc32_fifo_data_out[3] ;
    output \dc32_fifo_data_out[4] ;
    output \dc32_fifo_data_out[5] ;
    output \dc32_fifo_data_out[6] ;
    output \dc32_fifo_data_out[7] ;
    output \dc32_fifo_data_out[8] ;
    output \dc32_fifo_data_out[9] ;
    output \dc32_fifo_data_out[10] ;
    output \dc32_fifo_data_out[11] ;
    output \dc32_fifo_data_out[12] ;
    output \dc32_fifo_data_out[13] ;
    output \dc32_fifo_data_out[14] ;
    output \dc32_fifo_data_out[15] ;
    output \dc32_fifo_data_out[16] ;
    output \dc32_fifo_data_out[17] ;
    output \dc32_fifo_data_out[18] ;
    output \dc32_fifo_data_out[19] ;
    output \dc32_fifo_data_out[20] ;
    output \dc32_fifo_data_out[21] ;
    output \dc32_fifo_data_out[22] ;
    output \dc32_fifo_data_out[23] ;
    output \dc32_fifo_data_out[24] ;
    output \dc32_fifo_data_out[25] ;
    output \dc32_fifo_data_out[26] ;
    output \dc32_fifo_data_out[27] ;
    output \dc32_fifo_data_out[28] ;
    output \dc32_fifo_data_out[29] ;
    output \dc32_fifo_data_out[30] ;
    output \dc32_fifo_data_out[31] ;
    output n7_adj_6;
    output n8;
    input n25;
    input n5981;
    output \REG.mem_11_31 ;
    output \REG.mem_1_23 ;
    input n5980;
    output \REG.mem_11_30 ;
    output \REG.mem_6_6 ;
    output \REG.mem_7_6 ;
    output \REG.mem_5_6 ;
    output \REG.mem_4_6 ;
    input n5979;
    output \REG.mem_11_29 ;
    output \REG.mem_10_29 ;
    input n5978;
    input n5977;
    output \REG.mem_11_27 ;
    input n5976;
    output \REG.mem_11_26 ;
    input n5975;
    output \REG.mem_11_25 ;
    input n5974;
    output \REG.mem_11_24 ;
    output \REG.mem_9_29 ;
    output \REG.mem_8_29 ;
    input n5973;
    input n5972;
    output \REG.mem_11_22 ;
    output n29;
    output \REG.mem_8_17 ;
    output \REG.mem_9_17 ;
    output \REG.mem_10_17 ;
    output \REG.mem_11_17 ;
    output \REG.mem_1_24 ;
    input n5971;
    input n5970;
    output \REG.mem_11_20 ;
    output \REG.mem_6_31 ;
    output \REG.mem_7_31 ;
    output \REG.mem_5_31 ;
    output \REG.mem_4_31 ;
    output \wr_grey_sync_r[1] ;
    output n24;
    output n13;
    output n8_adj_7;
    output \REG.mem_6_23 ;
    output \REG.mem_7_23 ;
    output \REG.mem_5_23 ;
    output \REG.mem_4_23 ;
    output \REG.mem_10_6 ;
    output \REG.mem_11_6 ;
    input n5969;
    output \REG.mem_9_6 ;
    output \REG.mem_8_6 ;
    output \wr_grey_sync_r[2] ;
    output \wr_grey_sync_r[3] ;
    output \wr_grey_sync_r[4] ;
    input n5968;
    output \REG.mem_11_18 ;
    input n5967;
    input n5966;
    output \REG.mem_11_16 ;
    input n5965;
    input n5964;
    output \REG.mem_11_14 ;
    input n5963;
    input n5962;
    output \REG.mem_11_12 ;
    input n5961;
    input n5960;
    output \REG.mem_11_10 ;
    input n5959;
    output \REG.mem_11_9 ;
    input n5958;
    input n5957;
    output \REG.mem_11_7 ;
    input n5956;
    input n5955;
    output \REG.mem_11_5 ;
    input n5954;
    output \REG.mem_11_4 ;
    input n5953;
    output \REG.mem_11_3 ;
    output \REG.mem_10_22 ;
    input n5952;
    input n5951;
    output \REG.mem_11_1 ;
    input n5950;
    output \REG.mem_11_0 ;
    input n5949;
    output \REG.mem_10_31 ;
    input n5948;
    output \REG.mem_10_30 ;
    input n5947;
    input n5946;
    input n5945;
    output \REG.mem_10_27 ;
    output \REG.mem_9_22 ;
    output \REG.mem_8_22 ;
    input n5944;
    output \REG.mem_10_26 ;
    output \REG.mem_1_18 ;
    input n5943;
    output \REG.mem_10_25 ;
    input n5942;
    output \REG.mem_10_24 ;
    input n5611;
    output \REG.mem_6_24 ;
    output \REG.mem_7_24 ;
    output \REG.mem_5_24 ;
    output \REG.mem_4_24 ;
    output \REG.mem_1_4 ;
    output \REG.mem_9_24 ;
    output \REG.mem_8_24 ;
    output \REG.mem_6_0 ;
    output \REG.mem_7_0 ;
    output \REG.mem_5_0 ;
    output \REG.mem_4_0 ;
    output \REG.mem_10_4 ;
    input n5610;
    input n5941;
    input n5940;
    input n5939;
    input n5938;
    output \REG.mem_10_20 ;
    input n5937;
    input n5608;
    input n5604;
    input n5603;
    input n5602;
    input n5936;
    output \REG.mem_10_18 ;
    input n5935;
    input n5934;
    output \REG.mem_10_16 ;
    input n5933;
    output \REG.mem_1_17 ;
    output \REG.mem_9_4 ;
    output \REG.mem_8_4 ;
    output \REG.mem_6_17 ;
    output \REG.mem_7_17 ;
    output \REG.mem_4_17 ;
    output \REG.mem_5_17 ;
    input dc32_fifo_read_enable;
    input n5932;
    output \REG.mem_10_14 ;
    input n5931;
    input n5930;
    output \REG.mem_10_12 ;
    input n5929;
    input n5928;
    output \REG.mem_10_10 ;
    input n5927;
    output \REG.mem_10_9 ;
    input n5926;
    input n5925;
    output \REG.mem_10_7 ;
    input n5924;
    input n5923;
    output \REG.mem_10_5 ;
    input n5922;
    input n5921;
    output \REG.mem_10_3 ;
    input n5920;
    input n5919;
    output \REG.mem_10_1 ;
    input n5918;
    output \REG.mem_10_0 ;
    input n5917;
    output \REG.mem_9_31 ;
    input n5916;
    output \REG.mem_9_30 ;
    input n5915;
    input n5914;
    input n5913;
    output \REG.mem_9_27 ;
    input n5912;
    output \REG.mem_9_26 ;
    input n5911;
    output \REG.mem_9_25 ;
    input n5910;
    input n5909;
    input n5908;
    input n5907;
    input n5906;
    output \REG.mem_9_20 ;
    input n5905;
    input n5904;
    output \REG.mem_9_18 ;
    input n5903;
    input n5902;
    output \REG.mem_9_16 ;
    input n5901;
    input n5900;
    output \REG.mem_9_14 ;
    input n5899;
    input n5898;
    output \REG.mem_9_12 ;
    input n5897;
    input n5896;
    output \REG.mem_9_10 ;
    input n5895;
    output \REG.mem_9_9 ;
    input n5894;
    input n5893;
    output \REG.mem_9_7 ;
    input n5892;
    input n5891;
    input n5890;
    input n5889;
    output \REG.mem_9_3 ;
    input n5888;
    input n5887;
    output \REG.mem_9_1 ;
    input n5886;
    output \REG.mem_9_0 ;
    input n5885;
    output \REG.mem_8_31 ;
    input n5884;
    output \REG.mem_8_30 ;
    input n5883;
    input n5882;
    input n5881;
    output \REG.mem_8_27 ;
    input n5880;
    output \REG.mem_8_26 ;
    input n5879;
    output \REG.mem_8_25 ;
    input n5878;
    input n5877;
    input n5876;
    input n5875;
    input n5874;
    output \REG.mem_8_20 ;
    input n5873;
    input n5872;
    output \REG.mem_8_18 ;
    input n5871;
    input n5870;
    output \REG.mem_8_16 ;
    input n5869;
    input n5868;
    output \REG.mem_8_14 ;
    input n5867;
    input n5866;
    output \REG.mem_8_12 ;
    input n5865;
    input n5864;
    output \REG.mem_8_10 ;
    input n5863;
    output \REG.mem_8_9 ;
    input n5862;
    input n5861;
    output \REG.mem_8_7 ;
    input n5860;
    input n5859;
    input n5858;
    input n5857;
    output \REG.mem_8_3 ;
    input n5856;
    input n5855;
    output \REG.mem_8_1 ;
    input n5854;
    output \REG.mem_8_0 ;
    input n5853;
    input n5852;
    input n5851;
    output \REG.mem_7_29 ;
    input n5850;
    input n5849;
    input n5848;
    output \REG.mem_7_26 ;
    input n5847;
    output \REG.mem_7_25 ;
    input n5846;
    input n5845;
    input n5844;
    input n5843;
    input n5842;
    output \REG.mem_7_20 ;
    input n5841;
    input n5840;
    input n5839;
    input n5838;
    input n5837;
    output \REG.mem_7_15 ;
    input n5836;
    output \REG.mem_7_14 ;
    input n5835;
    input n5834;
    output \REG.mem_7_12 ;
    input n5833;
    output \REG.mem_7_11 ;
    input n5832;
    input n5831;
    input n5830;
    output \REG.mem_7_8 ;
    input n5829;
    input n5828;
    input n5827;
    output \REG.mem_7_5 ;
    input n5826;
    input n5825;
    output \REG.mem_7_3 ;
    input n5824;
    input n5823;
    input n5822;
    input n5821;
    input n5820;
    input n5819;
    output \REG.mem_6_29 ;
    input n5818;
    input n5817;
    input n5816;
    output \REG.mem_6_26 ;
    input n5815;
    output \REG.mem_6_25 ;
    input n5814;
    input n5813;
    input n5812;
    input n5811;
    input n5810;
    output \REG.mem_6_20 ;
    input n5809;
    input n5808;
    input n5807;
    input n5806;
    input n5805;
    output \REG.mem_6_15 ;
    input n5804;
    output \REG.mem_6_14 ;
    input n5803;
    input n5802;
    output \REG.mem_6_12 ;
    input n5801;
    output \REG.mem_6_11 ;
    input n5800;
    input n5799;
    input n5798;
    output \REG.mem_6_8 ;
    input n5797;
    input n5796;
    input n5795;
    output \REG.mem_6_5 ;
    input n5794;
    input n5793;
    output \REG.mem_6_3 ;
    input n5792;
    input n5791;
    input n5790;
    input n5789;
    input n5788;
    input n5600;
    output \REG.mem_1_3 ;
    input n5787;
    output \REG.mem_5_29 ;
    output n25_adj_8;
    output n9;
    input n5786;
    input n5785;
    input n5784;
    output \REG.mem_5_26 ;
    input n5783;
    output \REG.mem_5_25 ;
    input n5782;
    output \REG.mem_1_16 ;
    input n5781;
    input n5780;
    input n5779;
    input n5778;
    output \REG.mem_5_20 ;
    input n5777;
    input n5776;
    input n5775;
    input n5774;
    input n5773;
    output \REG.mem_5_15 ;
    input n5772;
    output \REG.mem_5_14 ;
    input n5771;
    input n5770;
    output \REG.mem_5_12 ;
    input n5769;
    output \REG.mem_5_11 ;
    output \REG.mem_1_25 ;
    input n5768;
    input n5767;
    input n5766;
    output \REG.mem_5_8 ;
    input n5765;
    output n10;
    output n26;
    input n5596;
    input n5764;
    input n5595;
    output \REG.mem_1_5 ;
    input n5594;
    input n5593;
    input n5590;
    input n5589;
    input n5588;
    input n5587;
    input n5763;
    output \REG.mem_5_5 ;
    output \REG.mem_4_26 ;
    input n5762;
    input n5761;
    output \REG.mem_5_3 ;
    input n5760;
    input n5759;
    input n5586;
    input n5758;
    input n5757;
    input n5756;
    input n5755;
    output \REG.mem_4_29 ;
    output \wr_addr_nxt_c[4] ;
    input n5754;
    input n5753;
    input n5752;
    input n5751;
    output \REG.mem_4_25 ;
    input n5750;
    input n5749;
    input n5748;
    input n5747;
    input n5585;
    output \REG.mem_1_29 ;
    input n5583;
    input n5582;
    input n5581;
    output \REG.mem_1_8 ;
    input n5580;
    input n5577;
    input n5746;
    output \REG.mem_4_20 ;
    input n5745;
    input n5744;
    input n5743;
    input n5742;
    input n5741;
    output \REG.mem_4_15 ;
    input n5740;
    output \REG.mem_4_14 ;
    input n5739;
    input n5738;
    output \REG.mem_4_12 ;
    input n5574;
    input n5572;
    input n5571;
    output \REG.mem_1_11 ;
    input n5737;
    output \REG.mem_4_11 ;
    input n5736;
    input n5735;
    input n5734;
    output \REG.mem_4_8 ;
    input n5733;
    input n5732;
    input n5731;
    output \REG.mem_4_5 ;
    input n5730;
    input n5729;
    output \REG.mem_4_3 ;
    input n5567;
    input n5565;
    output \REG.mem_1_20 ;
    input n5564;
    output \REG.mem_1_12 ;
    input n5560;
    input n5559;
    output \REG.mem_1_14 ;
    input n5558;
    output \REG.mem_1_15 ;
    input n5557;
    input n5556;
    input n5555;
    input n5554;
    input n5551;
    input n5550;
    input n5728;
    input n5727;
    input n5726;
    output n11;
    output n27;
    
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1 lscc_fifo_dc_inst (.dc32_fifo_data_in({dc32_fifo_data_in}), 
            .\REG.mem_1_9 (\REG.mem_1_9 ), .GND_net(GND_net), .\REG.mem_6_9 (\REG.mem_6_9 ), 
            .\REG.mem_7_9 (\REG.mem_7_9 ), .\REG.mem_4_9 (\REG.mem_4_9 ), 
            .\REG.mem_5_9 (\REG.mem_5_9 ), .\REG.mem_24_9 (\REG.mem_24_9 ), 
            .\REG.mem_25_9 (\REG.mem_25_9 ), .\REG.mem_1_31 (\REG.mem_1_31 ), 
            .\REG.mem_9_5 (\REG.mem_9_5 ), .\REG.mem_8_5 (\REG.mem_8_5 ), 
            .\REG.mem_26_9 (\REG.mem_26_9 ), .\REG.mem_27_9 (\REG.mem_27_9 ), 
            .rd_grey_sync_r({rd_grey_sync_r}), .\REG.mem_17_25 (\REG.mem_17_25 ), 
            .\REG.mem_6_16 (\REG.mem_6_16 ), .\REG.mem_7_16 (\REG.mem_7_16 ), 
            .\REG.mem_1_7 (\REG.mem_1_7 ), .\REG.mem_6_7 (\REG.mem_6_7 ), 
            .\REG.mem_7_7 (\REG.mem_7_7 ), .\REG.mem_4_7 (\REG.mem_4_7 ), 
            .\REG.mem_5_7 (\REG.mem_5_7 ), .\REG.mem_10_23 (\REG.mem_10_23 ), 
            .\REG.mem_11_23 (\REG.mem_11_23 ), .\REG.mem_5_16 (\REG.mem_5_16 ), 
            .\REG.mem_4_16 (\REG.mem_4_16 ), .\REG.mem_17_7 (\REG.mem_17_7 ), 
            .\REG.mem_22_7 (\REG.mem_22_7 ), .\REG.mem_23_7 (\REG.mem_23_7 ), 
            .\REG.mem_20_7 (\REG.mem_20_7 ), .\REG.mem_21_7 (\REG.mem_21_7 ), 
            .\REG.mem_9_23 (\REG.mem_9_23 ), .\REG.mem_8_23 (\REG.mem_8_23 ), 
            .n7(n7), .n23(n23), .FIFO_CLK_c(FIFO_CLK_c), .DEBUG_1_c(DEBUG_1_c), 
            .reset_per_frame(reset_per_frame), .wr_fifo_en_w(wr_fifo_en_w), 
            .\wr_addr_r[0] (\wr_addr_r[0] ), .\REG.mem_22_29 (\REG.mem_22_29 ), 
            .\REG.mem_23_29 (\REG.mem_23_29 ), .\REG.mem_21_29 (\REG.mem_21_29 ), 
            .\REG.mem_20_29 (\REG.mem_20_29 ), .DEBUG_5_c_0(DEBUG_5_c_0), 
            .SLM_CLK_c(SLM_CLK_c), .\REG.mem_26_21 (\REG.mem_26_21 ), .\REG.mem_27_21 (\REG.mem_27_21 ), 
            .\REG.mem_26_25 (\REG.mem_26_25 ), .\REG.mem_27_25 (\REG.mem_27_25 ), 
            .\REG.mem_25_25 (\REG.mem_25_25 ), .\REG.mem_24_25 (\REG.mem_24_25 ), 
            .\REG.mem_25_21 (\REG.mem_25_21 ), .\REG.mem_24_21 (\REG.mem_24_21 ), 
            .\REG.mem_1_10 (\REG.mem_1_10 ), .\REG.mem_6_10 (\REG.mem_6_10 ), 
            .\REG.mem_7_10 (\REG.mem_7_10 ), .\REG.mem_4_10 (\REG.mem_4_10 ), 
            .\REG.mem_5_10 (\REG.mem_5_10 ), .\REG.mem_1_26 (\REG.mem_1_26 ), 
            .n28(n28), .n12(n12), .dc32_fifo_empty(dc32_fifo_empty), .\wr_grey_sync_r[0] (\wr_grey_sync_r[0] ), 
            .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .dc32_fifo_almost_empty(dc32_fifo_almost_empty), .n32(n32), 
            .n16(n16), .\REG.mem_17_10 (\REG.mem_17_10 ), .\REG.mem_22_10 (\REG.mem_22_10 ), 
            .\REG.mem_23_10 (\REG.mem_23_10 ), .\REG.mem_20_10 (\REG.mem_20_10 ), 
            .\REG.mem_21_10 (\REG.mem_21_10 ), .dc32_fifo_full(dc32_fifo_full), 
            .\REG.mem_10_28 (\REG.mem_10_28 ), .\REG.mem_11_28 (\REG.mem_11_28 ), 
            .\REG.mem_9_28 (\REG.mem_9_28 ), .\REG.mem_8_28 (\REG.mem_8_28 ), 
            .\REG.mem_17_29 (\REG.mem_17_29 ), .\rd_addr_nxt_c_5__N_573[3] (\rd_addr_nxt_c_5__N_573[3] ), 
            .\rd_addr_nxt_c_5__N_573[1] (\rd_addr_nxt_c_5__N_573[1] ), .n6(n6), 
            .n22(n22), .\REG.mem_1_28 (\REG.mem_1_28 ), .\REG.mem_6_28 (\REG.mem_6_28 ), 
            .\REG.mem_7_28 (\REG.mem_7_28 ), .\REG.mem_4_28 (\REG.mem_4_28 ), 
            .\REG.mem_5_28 (\REG.mem_5_28 ), .\REG.mem_1_2 (\REG.mem_1_2 ), 
            .\REG.mem_6_2 (\REG.mem_6_2 ), .\REG.mem_7_2 (\REG.mem_7_2 ), 
            .\REG.mem_4_2 (\REG.mem_4_2 ), .\REG.mem_5_2 (\REG.mem_5_2 ), 
            .\REG.mem_1_22 (\REG.mem_1_22 ), .\REG.mem_6_22 (\REG.mem_6_22 ), 
            .\REG.mem_7_22 (\REG.mem_7_22 ), .\REG.mem_4_22 (\REG.mem_4_22 ), 
            .\REG.mem_5_22 (\REG.mem_5_22 ), .\REG.mem_17_22 (\REG.mem_17_22 ), 
            .\REG.mem_22_22 (\REG.mem_22_22 ), .\REG.mem_23_22 (\REG.mem_23_22 ), 
            .\REG.mem_20_22 (\REG.mem_20_22 ), .\REG.mem_21_22 (\REG.mem_21_22 ), 
            .\rd_addr_nxt_c_5__N_573[4] (\rd_addr_nxt_c_5__N_573[4] ), .\REG.mem_5_18 (\REG.mem_5_18 ), 
            .\REG.mem_4_18 (\REG.mem_4_18 ), .\REG.mem_6_4 (\REG.mem_6_4 ), 
            .\REG.mem_7_4 (\REG.mem_7_4 ), .\REG.mem_6_18 (\REG.mem_6_18 ), 
            .\REG.mem_7_18 (\REG.mem_7_18 ), .\REG.mem_10_8 (\REG.mem_10_8 ), 
            .\REG.mem_11_8 (\REG.mem_11_8 ), .\REG.mem_9_8 (\REG.mem_9_8 ), 
            .\REG.mem_8_8 (\REG.mem_8_8 ), .\REG.mem_5_4 (\REG.mem_5_4 ), 
            .\REG.mem_4_4 (\REG.mem_4_4 ), .\REG.mem_1_21 (\REG.mem_1_21 ), 
            .n7013(n7013), .n7012(n7012), .n7011(n7011), .n7010(n7010), 
            .n7009(n7009), .n7008(n7008), .wp_sync1_r({wp_sync1_r}), .n7007(n7007), 
            .n7006(n7006), .n7005(n7005), .n7004(n7004), .n7003(n7003), 
            .n7002(n7002), .n7000(n7000), .n6998(n6998), .n6997(n6997), 
            .n6996(n6996), .n6995(n6995), .n6994(n6994), .n6993(n6993), 
            .rp_sync1_r({rp_sync1_r}), .n6992(n6992), .n6991(n6991), .n6990(n6990), 
            .n6989(n6989), .\REG.mem_1_13 (\REG.mem_1_13 ), .n6930(n6930), 
            .n6928(n6928), .\wr_addr_r[5] (\wr_addr_r[5] ), .\REG.mem_6_30 (\REG.mem_6_30 ), 
            .\REG.mem_7_30 (\REG.mem_7_30 ), .n6493(n6493), .\REG.mem_27_31 (\REG.mem_27_31 ), 
            .n6492(n6492), .\REG.mem_27_30 (\REG.mem_27_30 ), .n6491(n6491), 
            .\REG.mem_27_29 (\REG.mem_27_29 ), .n6490(n6490), .\REG.mem_27_28 (\REG.mem_27_28 ), 
            .n6489(n6489), .\REG.mem_27_27 (\REG.mem_27_27 ), .n6488(n6488), 
            .\REG.mem_27_26 (\REG.mem_27_26 ), .n6487(n6487), .n6486(n6486), 
            .\REG.mem_27_24 (\REG.mem_27_24 ), .n6485(n6485), .\REG.mem_27_23 (\REG.mem_27_23 ), 
            .n6484(n6484), .\REG.mem_27_22 (\REG.mem_27_22 ), .n6483(n6483), 
            .n6482(n6482), .\REG.mem_27_20 (\REG.mem_27_20 ), .n6481(n6481), 
            .\REG.mem_27_19 (\REG.mem_27_19 ), .n6480(n6480), .\REG.mem_27_18 (\REG.mem_27_18 ), 
            .n6479(n6479), .\REG.mem_27_17 (\REG.mem_27_17 ), .n6478(n6478), 
            .\REG.mem_27_16 (\REG.mem_27_16 ), .n6477(n6477), .\REG.mem_27_15 (\REG.mem_27_15 ), 
            .n6476(n6476), .\REG.mem_27_14 (\REG.mem_27_14 ), .n6475(n6475), 
            .\REG.mem_27_13 (\REG.mem_27_13 ), .n6474(n6474), .\REG.mem_27_12 (\REG.mem_27_12 ), 
            .n6473(n6473), .\REG.mem_27_11 (\REG.mem_27_11 ), .n6472(n6472), 
            .\REG.mem_27_10 (\REG.mem_27_10 ), .n6471(n6471), .n6470(n6470), 
            .\REG.mem_27_8 (\REG.mem_27_8 ), .n6469(n6469), .\REG.mem_27_7 (\REG.mem_27_7 ), 
            .n6468(n6468), .\REG.mem_27_6 (\REG.mem_27_6 ), .n6467(n6467), 
            .\REG.mem_27_5 (\REG.mem_27_5 ), .n6466(n6466), .\REG.mem_27_4 (\REG.mem_27_4 ), 
            .n6465(n6465), .\REG.mem_27_3 (\REG.mem_27_3 ), .n6464(n6464), 
            .\REG.mem_27_2 (\REG.mem_27_2 ), .n6463(n6463), .\REG.mem_27_1 (\REG.mem_27_1 ), 
            .n6462(n6462), .\REG.mem_27_0 (\REG.mem_27_0 ), .n6461(n6461), 
            .\REG.mem_26_31 (\REG.mem_26_31 ), .n6460(n6460), .\REG.mem_26_30 (\REG.mem_26_30 ), 
            .n6459(n6459), .\REG.mem_26_29 (\REG.mem_26_29 ), .n6458(n6458), 
            .\REG.mem_26_28 (\REG.mem_26_28 ), .n6457(n6457), .\REG.mem_26_27 (\REG.mem_26_27 ), 
            .n6456(n6456), .\REG.mem_26_26 (\REG.mem_26_26 ), .n6455(n6455), 
            .n6454(n6454), .\REG.mem_26_24 (\REG.mem_26_24 ), .n6453(n6453), 
            .\REG.mem_26_23 (\REG.mem_26_23 ), .n6452(n6452), .\REG.mem_26_22 (\REG.mem_26_22 ), 
            .n6451(n6451), .n6450(n6450), .\REG.mem_26_20 (\REG.mem_26_20 ), 
            .n6449(n6449), .\REG.mem_26_19 (\REG.mem_26_19 ), .n6448(n6448), 
            .\REG.mem_26_18 (\REG.mem_26_18 ), .n6447(n6447), .\REG.mem_26_17 (\REG.mem_26_17 ), 
            .n6446(n6446), .\REG.mem_26_16 (\REG.mem_26_16 ), .n6445(n6445), 
            .\REG.mem_26_15 (\REG.mem_26_15 ), .n6444(n6444), .\REG.mem_26_14 (\REG.mem_26_14 ), 
            .n6443(n6443), .\REG.mem_26_13 (\REG.mem_26_13 ), .n6442(n6442), 
            .\REG.mem_26_12 (\REG.mem_26_12 ), .n6441(n6441), .\REG.mem_26_11 (\REG.mem_26_11 ), 
            .n6440(n6440), .\REG.mem_26_10 (\REG.mem_26_10 ), .n6439(n6439), 
            .n6438(n6438), .\REG.mem_26_8 (\REG.mem_26_8 ), .n6437(n6437), 
            .\REG.mem_26_7 (\REG.mem_26_7 ), .n6436(n6436), .\REG.mem_26_6 (\REG.mem_26_6 ), 
            .n6435(n6435), .\REG.mem_26_5 (\REG.mem_26_5 ), .n6434(n6434), 
            .\REG.mem_26_4 (\REG.mem_26_4 ), .n6433(n6433), .\REG.mem_26_3 (\REG.mem_26_3 ), 
            .n6432(n6432), .\REG.mem_26_2 (\REG.mem_26_2 ), .n6431(n6431), 
            .\REG.mem_26_1 (\REG.mem_26_1 ), .n6430(n6430), .\REG.mem_26_0 (\REG.mem_26_0 ), 
            .n6429(n6429), .\REG.mem_25_31 (\REG.mem_25_31 ), .n6428(n6428), 
            .\REG.mem_25_30 (\REG.mem_25_30 ), .n6427(n6427), .\REG.mem_25_29 (\REG.mem_25_29 ), 
            .n6426(n6426), .\REG.mem_25_28 (\REG.mem_25_28 ), .n6425(n6425), 
            .\REG.mem_25_27 (\REG.mem_25_27 ), .n6424(n6424), .\REG.mem_25_26 (\REG.mem_25_26 ), 
            .n6423(n6423), .n6422(n6422), .\REG.mem_25_24 (\REG.mem_25_24 ), 
            .n6421(n6421), .\REG.mem_25_23 (\REG.mem_25_23 ), .n6420(n6420), 
            .\REG.mem_25_22 (\REG.mem_25_22 ), .n6419(n6419), .n6418(n6418), 
            .\REG.mem_25_20 (\REG.mem_25_20 ), .n6417(n6417), .\REG.mem_25_19 (\REG.mem_25_19 ), 
            .n6416(n6416), .\REG.mem_25_18 (\REG.mem_25_18 ), .n6415(n6415), 
            .\REG.mem_25_17 (\REG.mem_25_17 ), .n6414(n6414), .\REG.mem_25_16 (\REG.mem_25_16 ), 
            .n6413(n6413), .\REG.mem_25_15 (\REG.mem_25_15 ), .n6412(n6412), 
            .\REG.mem_25_14 (\REG.mem_25_14 ), .n6411(n6411), .\REG.mem_25_13 (\REG.mem_25_13 ), 
            .n6410(n6410), .\REG.mem_25_12 (\REG.mem_25_12 ), .n6409(n6409), 
            .\REG.mem_25_11 (\REG.mem_25_11 ), .n6408(n6408), .\REG.mem_25_10 (\REG.mem_25_10 ), 
            .n6407(n6407), .n6406(n6406), .\REG.mem_25_8 (\REG.mem_25_8 ), 
            .n6405(n6405), .\REG.mem_25_7 (\REG.mem_25_7 ), .n6404(n6404), 
            .\REG.mem_25_6 (\REG.mem_25_6 ), .n6403(n6403), .\REG.mem_25_5 (\REG.mem_25_5 ), 
            .n6402(n6402), .\REG.mem_25_4 (\REG.mem_25_4 ), .n6401(n6401), 
            .\REG.mem_25_3 (\REG.mem_25_3 ), .n6400(n6400), .\REG.mem_25_2 (\REG.mem_25_2 ), 
            .n6399(n6399), .\REG.mem_25_1 (\REG.mem_25_1 ), .n6398(n6398), 
            .\REG.mem_25_0 (\REG.mem_25_0 ), .n6397(n6397), .\REG.mem_24_31 (\REG.mem_24_31 ), 
            .n6396(n6396), .\REG.mem_24_30 (\REG.mem_24_30 ), .n6395(n6395), 
            .\REG.mem_24_29 (\REG.mem_24_29 ), .n6394(n6394), .\REG.mem_24_28 (\REG.mem_24_28 ), 
            .n6393(n6393), .\REG.mem_24_27 (\REG.mem_24_27 ), .n6392(n6392), 
            .\REG.mem_24_26 (\REG.mem_24_26 ), .n6391(n6391), .n6390(n6390), 
            .\REG.mem_24_24 (\REG.mem_24_24 ), .n6389(n6389), .\REG.mem_24_23 (\REG.mem_24_23 ), 
            .n6388(n6388), .\REG.mem_24_22 (\REG.mem_24_22 ), .n6387(n6387), 
            .n6386(n6386), .\REG.mem_24_20 (\REG.mem_24_20 ), .n6385(n6385), 
            .\REG.mem_24_19 (\REG.mem_24_19 ), .n6384(n6384), .\REG.mem_24_18 (\REG.mem_24_18 ), 
            .n6383(n6383), .\REG.mem_24_17 (\REG.mem_24_17 ), .n6382(n6382), 
            .\REG.mem_24_16 (\REG.mem_24_16 ), .n6381(n6381), .\REG.mem_24_15 (\REG.mem_24_15 ), 
            .n6380(n6380), .\REG.mem_24_14 (\REG.mem_24_14 ), .n6379(n6379), 
            .\REG.mem_24_13 (\REG.mem_24_13 ), .n6378(n6378), .\REG.mem_24_12 (\REG.mem_24_12 ), 
            .n6377(n6377), .\REG.mem_24_11 (\REG.mem_24_11 ), .n6376(n6376), 
            .\REG.mem_24_10 (\REG.mem_24_10 ), .n6375(n6375), .n6374(n6374), 
            .\REG.mem_24_8 (\REG.mem_24_8 ), .n6373(n6373), .\REG.mem_24_7 (\REG.mem_24_7 ), 
            .n6372(n6372), .\REG.mem_24_6 (\REG.mem_24_6 ), .n6371(n6371), 
            .\REG.mem_24_5 (\REG.mem_24_5 ), .n6370(n6370), .\REG.mem_24_4 (\REG.mem_24_4 ), 
            .n6369(n6369), .\REG.mem_24_3 (\REG.mem_24_3 ), .n6368(n6368), 
            .\REG.mem_24_2 (\REG.mem_24_2 ), .n6367(n6367), .\REG.mem_24_1 (\REG.mem_24_1 ), 
            .n6366(n6366), .\REG.mem_24_0 (\REG.mem_24_0 ), .n6365(n6365), 
            .\REG.mem_23_31 (\REG.mem_23_31 ), .n6364(n6364), .\REG.mem_23_30 (\REG.mem_23_30 ), 
            .n6363(n6363), .n6362(n6362), .\REG.mem_23_28 (\REG.mem_23_28 ), 
            .n6361(n6361), .\REG.mem_23_27 (\REG.mem_23_27 ), .n6360(n6360), 
            .\REG.mem_23_26 (\REG.mem_23_26 ), .n6359(n6359), .\REG.mem_23_25 (\REG.mem_23_25 ), 
            .n6358(n6358), .\REG.mem_23_24 (\REG.mem_23_24 ), .n6357(n6357), 
            .\REG.mem_23_23 (\REG.mem_23_23 ), .n6356(n6356), .n6355(n6355), 
            .\REG.mem_23_21 (\REG.mem_23_21 ), .n6354(n6354), .\REG.mem_23_20 (\REG.mem_23_20 ), 
            .n6353(n6353), .\REG.mem_23_19 (\REG.mem_23_19 ), .n6352(n6352), 
            .\REG.mem_23_18 (\REG.mem_23_18 ), .n6351(n6351), .\REG.mem_23_17 (\REG.mem_23_17 ), 
            .n6350(n6350), .\REG.mem_23_16 (\REG.mem_23_16 ), .n6349(n6349), 
            .\REG.mem_23_15 (\REG.mem_23_15 ), .n6348(n6348), .\REG.mem_23_14 (\REG.mem_23_14 ), 
            .n6347(n6347), .\REG.mem_23_13 (\REG.mem_23_13 ), .n6346(n6346), 
            .\REG.mem_23_12 (\REG.mem_23_12 ), .n6345(n6345), .\REG.mem_23_11 (\REG.mem_23_11 ), 
            .n6344(n6344), .n6343(n6343), .\REG.mem_23_9 (\REG.mem_23_9 ), 
            .n6342(n6342), .\REG.mem_23_8 (\REG.mem_23_8 ), .n6341(n6341), 
            .n6340(n6340), .\REG.mem_23_6 (\REG.mem_23_6 ), .n6339(n6339), 
            .\REG.mem_23_5 (\REG.mem_23_5 ), .n6338(n6338), .\REG.mem_23_4 (\REG.mem_23_4 ), 
            .n6337(n6337), .\REG.mem_23_3 (\REG.mem_23_3 ), .n6336(n6336), 
            .\REG.mem_23_2 (\REG.mem_23_2 ), .n6335(n6335), .\REG.mem_23_1 (\REG.mem_23_1 ), 
            .n6334(n6334), .\REG.mem_23_0 (\REG.mem_23_0 ), .n6333(n6333), 
            .\REG.mem_22_31 (\REG.mem_22_31 ), .n6332(n6332), .\REG.mem_22_30 (\REG.mem_22_30 ), 
            .n6331(n6331), .n6330(n6330), .\REG.mem_22_28 (\REG.mem_22_28 ), 
            .n6329(n6329), .\REG.mem_22_27 (\REG.mem_22_27 ), .n6328(n6328), 
            .\REG.mem_22_26 (\REG.mem_22_26 ), .n6327(n6327), .\REG.mem_22_25 (\REG.mem_22_25 ), 
            .n6326(n6326), .\REG.mem_22_24 (\REG.mem_22_24 ), .n6325(n6325), 
            .\REG.mem_22_23 (\REG.mem_22_23 ), .n6324(n6324), .n6323(n6323), 
            .\REG.mem_22_21 (\REG.mem_22_21 ), .n6322(n6322), .\REG.mem_22_20 (\REG.mem_22_20 ), 
            .n6321(n6321), .\REG.mem_22_19 (\REG.mem_22_19 ), .n6320(n6320), 
            .\REG.mem_22_18 (\REG.mem_22_18 ), .n6319(n6319), .\REG.mem_22_17 (\REG.mem_22_17 ), 
            .n6318(n6318), .\REG.mem_22_16 (\REG.mem_22_16 ), .n6317(n6317), 
            .\REG.mem_22_15 (\REG.mem_22_15 ), .n6316(n6316), .\REG.mem_22_14 (\REG.mem_22_14 ), 
            .n6315(n6315), .\REG.mem_22_13 (\REG.mem_22_13 ), .n6314(n6314), 
            .\REG.mem_22_12 (\REG.mem_22_12 ), .n6313(n6313), .\REG.mem_22_11 (\REG.mem_22_11 ), 
            .n6312(n6312), .n6311(n6311), .\REG.mem_22_9 (\REG.mem_22_9 ), 
            .n6310(n6310), .\REG.mem_22_8 (\REG.mem_22_8 ), .n6309(n6309), 
            .n6308(n6308), .\REG.mem_22_6 (\REG.mem_22_6 ), .n6307(n6307), 
            .\REG.mem_22_5 (\REG.mem_22_5 ), .n6306(n6306), .\REG.mem_22_4 (\REG.mem_22_4 ), 
            .n6305(n6305), .\REG.mem_22_3 (\REG.mem_22_3 ), .n6304(n6304), 
            .\REG.mem_22_2 (\REG.mem_22_2 ), .n6303(n6303), .\REG.mem_22_1 (\REG.mem_22_1 ), 
            .n6302(n6302), .\REG.mem_22_0 (\REG.mem_22_0 ), .n6301(n6301), 
            .\REG.mem_21_31 (\REG.mem_21_31 ), .n6300(n6300), .\REG.mem_21_30 (\REG.mem_21_30 ), 
            .n6299(n6299), .n6298(n6298), .\REG.mem_21_28 (\REG.mem_21_28 ), 
            .n6297(n6297), .\REG.mem_21_27 (\REG.mem_21_27 ), .n6296(n6296), 
            .\REG.mem_21_26 (\REG.mem_21_26 ), .n6295(n6295), .\REG.mem_21_25 (\REG.mem_21_25 ), 
            .n6294(n6294), .\REG.mem_21_24 (\REG.mem_21_24 ), .n6293(n6293), 
            .\REG.mem_21_23 (\REG.mem_21_23 ), .n6292(n6292), .n6291(n6291), 
            .\REG.mem_21_21 (\REG.mem_21_21 ), .n6290(n6290), .\REG.mem_21_20 (\REG.mem_21_20 ), 
            .n6289(n6289), .\REG.mem_21_19 (\REG.mem_21_19 ), .n6288(n6288), 
            .\REG.mem_21_18 (\REG.mem_21_18 ), .n6287(n6287), .\REG.mem_21_17 (\REG.mem_21_17 ), 
            .n6286(n6286), .\REG.mem_21_16 (\REG.mem_21_16 ), .n6285(n6285), 
            .\REG.mem_21_15 (\REG.mem_21_15 ), .n6284(n6284), .\REG.mem_21_14 (\REG.mem_21_14 ), 
            .n6283(n6283), .\REG.mem_21_13 (\REG.mem_21_13 ), .n6282(n6282), 
            .\REG.mem_21_12 (\REG.mem_21_12 ), .n6281(n6281), .\REG.mem_21_11 (\REG.mem_21_11 ), 
            .n6280(n6280), .n6279(n6279), .\REG.mem_21_9 (\REG.mem_21_9 ), 
            .n6278(n6278), .\REG.mem_21_8 (\REG.mem_21_8 ), .n6277(n6277), 
            .n6276(n6276), .\REG.mem_21_6 (\REG.mem_21_6 ), .n6275(n6275), 
            .\REG.mem_21_5 (\REG.mem_21_5 ), .n6274(n6274), .\REG.mem_21_4 (\REG.mem_21_4 ), 
            .n6273(n6273), .\REG.mem_21_3 (\REG.mem_21_3 ), .n6272(n6272), 
            .\REG.mem_21_2 (\REG.mem_21_2 ), .n6271(n6271), .\REG.mem_21_1 (\REG.mem_21_1 ), 
            .n6270(n6270), .\REG.mem_21_0 (\REG.mem_21_0 ), .n6269(n6269), 
            .\REG.mem_20_31 (\REG.mem_20_31 ), .n6268(n6268), .\REG.mem_20_30 (\REG.mem_20_30 ), 
            .n6267(n6267), .n6266(n6266), .\REG.mem_20_28 (\REG.mem_20_28 ), 
            .n6265(n6265), .\REG.mem_20_27 (\REG.mem_20_27 ), .n6264(n6264), 
            .\REG.mem_20_26 (\REG.mem_20_26 ), .n6263(n6263), .\REG.mem_20_25 (\REG.mem_20_25 ), 
            .n6262(n6262), .\REG.mem_20_24 (\REG.mem_20_24 ), .n6261(n6261), 
            .\REG.mem_20_23 (\REG.mem_20_23 ), .n6260(n6260), .n6259(n6259), 
            .\REG.mem_20_21 (\REG.mem_20_21 ), .n6258(n6258), .\REG.mem_20_20 (\REG.mem_20_20 ), 
            .n6257(n6257), .\REG.mem_20_19 (\REG.mem_20_19 ), .n6256(n6256), 
            .\REG.mem_20_18 (\REG.mem_20_18 ), .n6255(n6255), .\REG.mem_20_17 (\REG.mem_20_17 ), 
            .n6254(n6254), .\REG.mem_20_16 (\REG.mem_20_16 ), .n6253(n6253), 
            .\REG.mem_20_15 (\REG.mem_20_15 ), .n6252(n6252), .\REG.mem_20_14 (\REG.mem_20_14 ), 
            .n6251(n6251), .\REG.mem_20_13 (\REG.mem_20_13 ), .n6250(n6250), 
            .\REG.mem_20_12 (\REG.mem_20_12 ), .n6249(n6249), .\REG.mem_20_11 (\REG.mem_20_11 ), 
            .n6248(n6248), .n6247(n6247), .\REG.mem_20_9 (\REG.mem_20_9 ), 
            .n6246(n6246), .\REG.mem_20_8 (\REG.mem_20_8 ), .n6245(n6245), 
            .n6244(n6244), .\REG.mem_20_6 (\REG.mem_20_6 ), .n6243(n6243), 
            .\REG.mem_20_5 (\REG.mem_20_5 ), .n6242(n6242), .\REG.mem_20_4 (\REG.mem_20_4 ), 
            .n6241(n6241), .\REG.mem_20_3 (\REG.mem_20_3 ), .n6240(n6240), 
            .\REG.mem_20_2 (\REG.mem_20_2 ), .n6239(n6239), .\REG.mem_20_1 (\REG.mem_20_1 ), 
            .n6238(n6238), .\REG.mem_20_0 (\REG.mem_20_0 ), .n6173(n6173), 
            .\REG.mem_17_31 (\REG.mem_17_31 ), .n6172(n6172), .\REG.mem_17_30 (\REG.mem_17_30 ), 
            .n6171(n6171), .n6170(n6170), .\REG.mem_17_28 (\REG.mem_17_28 ), 
            .n6169(n6169), .\REG.mem_17_27 (\REG.mem_17_27 ), .n6168(n6168), 
            .\REG.mem_17_26 (\REG.mem_17_26 ), .n6167(n6167), .n6166(n6166), 
            .\REG.mem_17_24 (\REG.mem_17_24 ), .n6165(n6165), .\REG.mem_17_23 (\REG.mem_17_23 ), 
            .n6164(n6164), .n6163(n6163), .\REG.mem_17_21 (\REG.mem_17_21 ), 
            .n6162(n6162), .\REG.mem_17_20 (\REG.mem_17_20 ), .n6161(n6161), 
            .\REG.mem_17_19 (\REG.mem_17_19 ), .n6160(n6160), .\REG.mem_17_18 (\REG.mem_17_18 ), 
            .n6159(n6159), .\REG.mem_17_17 (\REG.mem_17_17 ), .n6158(n6158), 
            .\REG.mem_17_16 (\REG.mem_17_16 ), .n6157(n6157), .\REG.mem_17_15 (\REG.mem_17_15 ), 
            .n6156(n6156), .\REG.mem_17_14 (\REG.mem_17_14 ), .n6155(n6155), 
            .\REG.mem_17_13 (\REG.mem_17_13 ), .n6154(n6154), .\REG.mem_17_12 (\REG.mem_17_12 ), 
            .n6153(n6153), .\REG.mem_17_11 (\REG.mem_17_11 ), .n6152(n6152), 
            .n6151(n6151), .\REG.mem_17_9 (\REG.mem_17_9 ), .n6150(n6150), 
            .\REG.mem_17_8 (\REG.mem_17_8 ), .n6149(n6149), .n6148(n6148), 
            .\REG.mem_17_6 (\REG.mem_17_6 ), .n6147(n6147), .\REG.mem_17_5 (\REG.mem_17_5 ), 
            .n6146(n6146), .\REG.mem_17_4 (\REG.mem_17_4 ), .n6145(n6145), 
            .\REG.mem_17_3 (\REG.mem_17_3 ), .n6144(n6144), .\REG.mem_17_2 (\REG.mem_17_2 ), 
            .n6143(n6143), .\REG.mem_17_1 (\REG.mem_17_1 ), .n6142(n6142), 
            .\REG.mem_17_0 (\REG.mem_17_0 ), .\REG.mem_5_30 (\REG.mem_5_30 ), 
            .\REG.mem_4_30 (\REG.mem_4_30 ), .\REG.mem_1_1 (\REG.mem_1_1 ), 
            .\REG.mem_6_1 (\REG.mem_6_1 ), .\REG.mem_7_1 (\REG.mem_7_1 ), 
            .\REG.mem_4_1 (\REG.mem_4_1 ), .\REG.mem_5_1 (\REG.mem_5_1 ), 
            .\REG.mem_6_21 (\REG.mem_6_21 ), .\REG.mem_7_21 (\REG.mem_7_21 ), 
            .\REG.mem_5_21 (\REG.mem_5_21 ), .\REG.mem_4_21 (\REG.mem_4_21 ), 
            .\REG.mem_1_30 (\REG.mem_1_30 ), .\REG.mem_10_21 (\REG.mem_10_21 ), 
            .\REG.mem_11_21 (\REG.mem_11_21 ), .\REG.mem_1_19 (\REG.mem_1_19 ), 
            .\REG.mem_6_19 (\REG.mem_6_19 ), .\REG.mem_7_19 (\REG.mem_7_19 ), 
            .\REG.mem_5_19 (\REG.mem_5_19 ), .\REG.mem_4_19 (\REG.mem_4_19 ), 
            .\REG.mem_9_21 (\REG.mem_9_21 ), .\REG.mem_8_21 (\REG.mem_8_21 ), 
            .\wr_addr_p1_w[0] (\wr_addr_p1_w[0] ), .\REG.mem_6_13 (\REG.mem_6_13 ), 
            .\REG.mem_7_13 (\REG.mem_7_13 ), .\REG.mem_5_13 (\REG.mem_5_13 ), 
            .\REG.mem_4_13 (\REG.mem_4_13 ), .\REG.mem_10_13 (\REG.mem_10_13 ), 
            .\REG.mem_11_13 (\REG.mem_11_13 ), .\REG.mem_9_13 (\REG.mem_9_13 ), 
            .\REG.mem_8_13 (\REG.mem_8_13 ), .\REG.mem_10_19 (\REG.mem_10_19 ), 
            .\REG.mem_11_19 (\REG.mem_11_19 ), .\REG.mem_9_19 (\REG.mem_9_19 ), 
            .\REG.mem_8_19 (\REG.mem_8_19 ), .\REG.mem_1_27 (\REG.mem_1_27 ), 
            .\REG.mem_6_27 (\REG.mem_6_27 ), .\REG.mem_7_27 (\REG.mem_7_27 ), 
            .\REG.mem_4_27 (\REG.mem_4_27 ), .\REG.mem_5_27 (\REG.mem_5_27 ), 
            .\REG.mem_1_6 (\REG.mem_1_6 ), .\REG.mem_8_2 (\REG.mem_8_2 ), 
            .\REG.mem_9_2 (\REG.mem_9_2 ), .\REG.mem_10_2 (\REG.mem_10_2 ), 
            .\REG.mem_11_2 (\REG.mem_11_2 ), .\wr_addr_nxt_c[2] (\wr_addr_nxt_c[2] ), 
            .VCC_net(VCC_net), .dc32_fifo_write_enable(dc32_fifo_write_enable), 
            .\REG.mem_1_0 (\REG.mem_1_0 ), .\REG.mem_10_15 (\REG.mem_10_15 ), 
            .\REG.mem_11_15 (\REG.mem_11_15 ), .\REG.mem_9_15 (\REG.mem_9_15 ), 
            .\REG.mem_8_15 (\REG.mem_8_15 ), .\dc32_fifo_data_out[1] (\dc32_fifo_data_out[1] ), 
            .\REG.mem_10_11 (\REG.mem_10_11 ), .\REG.mem_11_11 (\REG.mem_11_11 ), 
            .\REG.mem_9_11 (\REG.mem_9_11 ), .\REG.mem_8_11 (\REG.mem_8_11 ), 
            .\dc32_fifo_data_out[2] (\dc32_fifo_data_out[2] ), .\dc32_fifo_data_out[3] (\dc32_fifo_data_out[3] ), 
            .\dc32_fifo_data_out[4] (\dc32_fifo_data_out[4] ), .\dc32_fifo_data_out[5] (\dc32_fifo_data_out[5] ), 
            .\dc32_fifo_data_out[6] (\dc32_fifo_data_out[6] ), .\dc32_fifo_data_out[7] (\dc32_fifo_data_out[7] ), 
            .\dc32_fifo_data_out[8] (\dc32_fifo_data_out[8] ), .\dc32_fifo_data_out[9] (\dc32_fifo_data_out[9] ), 
            .\dc32_fifo_data_out[10] (\dc32_fifo_data_out[10] ), .\dc32_fifo_data_out[11] (\dc32_fifo_data_out[11] ), 
            .\dc32_fifo_data_out[12] (\dc32_fifo_data_out[12] ), .\dc32_fifo_data_out[13] (\dc32_fifo_data_out[13] ), 
            .\dc32_fifo_data_out[14] (\dc32_fifo_data_out[14] ), .\dc32_fifo_data_out[15] (\dc32_fifo_data_out[15] ), 
            .\dc32_fifo_data_out[16] (\dc32_fifo_data_out[16] ), .\dc32_fifo_data_out[17] (\dc32_fifo_data_out[17] ), 
            .\dc32_fifo_data_out[18] (\dc32_fifo_data_out[18] ), .\dc32_fifo_data_out[19] (\dc32_fifo_data_out[19] ), 
            .\dc32_fifo_data_out[20] (\dc32_fifo_data_out[20] ), .\dc32_fifo_data_out[21] (\dc32_fifo_data_out[21] ), 
            .\dc32_fifo_data_out[22] (\dc32_fifo_data_out[22] ), .\dc32_fifo_data_out[23] (\dc32_fifo_data_out[23] ), 
            .\dc32_fifo_data_out[24] (\dc32_fifo_data_out[24] ), .\dc32_fifo_data_out[25] (\dc32_fifo_data_out[25] ), 
            .\dc32_fifo_data_out[26] (\dc32_fifo_data_out[26] ), .\dc32_fifo_data_out[27] (\dc32_fifo_data_out[27] ), 
            .\dc32_fifo_data_out[28] (\dc32_fifo_data_out[28] ), .\dc32_fifo_data_out[29] (\dc32_fifo_data_out[29] ), 
            .\dc32_fifo_data_out[30] (\dc32_fifo_data_out[30] ), .\dc32_fifo_data_out[31] (\dc32_fifo_data_out[31] ), 
            .n7_adj_3(n7_adj_6), .n8(n8), .n25(n25), .n5981(n5981), 
            .\REG.mem_11_31 (\REG.mem_11_31 ), .\REG.mem_1_23 (\REG.mem_1_23 ), 
            .n5980(n5980), .\REG.mem_11_30 (\REG.mem_11_30 ), .\REG.mem_6_6 (\REG.mem_6_6 ), 
            .\REG.mem_7_6 (\REG.mem_7_6 ), .\REG.mem_5_6 (\REG.mem_5_6 ), 
            .\REG.mem_4_6 (\REG.mem_4_6 ), .n5979(n5979), .\REG.mem_11_29 (\REG.mem_11_29 ), 
            .\REG.mem_10_29 (\REG.mem_10_29 ), .n5978(n5978), .n5977(n5977), 
            .\REG.mem_11_27 (\REG.mem_11_27 ), .n5976(n5976), .\REG.mem_11_26 (\REG.mem_11_26 ), 
            .n5975(n5975), .\REG.mem_11_25 (\REG.mem_11_25 ), .n5974(n5974), 
            .\REG.mem_11_24 (\REG.mem_11_24 ), .\REG.mem_9_29 (\REG.mem_9_29 ), 
            .\REG.mem_8_29 (\REG.mem_8_29 ), .n5973(n5973), .n5972(n5972), 
            .\REG.mem_11_22 (\REG.mem_11_22 ), .n29(n29), .\REG.mem_8_17 (\REG.mem_8_17 ), 
            .\REG.mem_9_17 (\REG.mem_9_17 ), .\REG.mem_10_17 (\REG.mem_10_17 ), 
            .\REG.mem_11_17 (\REG.mem_11_17 ), .\REG.mem_1_24 (\REG.mem_1_24 ), 
            .n5971(n5971), .n5970(n5970), .\REG.mem_11_20 (\REG.mem_11_20 ), 
            .\REG.mem_6_31 (\REG.mem_6_31 ), .\REG.mem_7_31 (\REG.mem_7_31 ), 
            .\REG.mem_5_31 (\REG.mem_5_31 ), .\REG.mem_4_31 (\REG.mem_4_31 ), 
            .\wr_grey_sync_r[1] (\wr_grey_sync_r[1] ), .n24(n24), .n13(n13), 
            .n8_adj_4(n8_adj_7), .\REG.mem_6_23 (\REG.mem_6_23 ), .\REG.mem_7_23 (\REG.mem_7_23 ), 
            .\REG.mem_5_23 (\REG.mem_5_23 ), .\REG.mem_4_23 (\REG.mem_4_23 ), 
            .\REG.mem_10_6 (\REG.mem_10_6 ), .\REG.mem_11_6 (\REG.mem_11_6 ), 
            .n5969(n5969), .\REG.mem_9_6 (\REG.mem_9_6 ), .\REG.mem_8_6 (\REG.mem_8_6 ), 
            .\wr_grey_sync_r[2] (\wr_grey_sync_r[2] ), .\wr_grey_sync_r[3] (\wr_grey_sync_r[3] ), 
            .\wr_grey_sync_r[4] (\wr_grey_sync_r[4] ), .n5968(n5968), .\REG.mem_11_18 (\REG.mem_11_18 ), 
            .n5967(n5967), .n5966(n5966), .\REG.mem_11_16 (\REG.mem_11_16 ), 
            .n5965(n5965), .n5964(n5964), .\REG.mem_11_14 (\REG.mem_11_14 ), 
            .n5963(n5963), .n5962(n5962), .\REG.mem_11_12 (\REG.mem_11_12 ), 
            .n5961(n5961), .n5960(n5960), .\REG.mem_11_10 (\REG.mem_11_10 ), 
            .n5959(n5959), .\REG.mem_11_9 (\REG.mem_11_9 ), .n5958(n5958), 
            .n5957(n5957), .\REG.mem_11_7 (\REG.mem_11_7 ), .n5956(n5956), 
            .n5955(n5955), .\REG.mem_11_5 (\REG.mem_11_5 ), .n5954(n5954), 
            .\REG.mem_11_4 (\REG.mem_11_4 ), .n5953(n5953), .\REG.mem_11_3 (\REG.mem_11_3 ), 
            .\REG.mem_10_22 (\REG.mem_10_22 ), .n5952(n5952), .n5951(n5951), 
            .\REG.mem_11_1 (\REG.mem_11_1 ), .n5950(n5950), .\REG.mem_11_0 (\REG.mem_11_0 ), 
            .n5949(n5949), .\REG.mem_10_31 (\REG.mem_10_31 ), .n5948(n5948), 
            .\REG.mem_10_30 (\REG.mem_10_30 ), .n5947(n5947), .n5946(n5946), 
            .n5945(n5945), .\REG.mem_10_27 (\REG.mem_10_27 ), .\REG.mem_9_22 (\REG.mem_9_22 ), 
            .\REG.mem_8_22 (\REG.mem_8_22 ), .n5944(n5944), .\REG.mem_10_26 (\REG.mem_10_26 ), 
            .\REG.mem_1_18 (\REG.mem_1_18 ), .n5943(n5943), .\REG.mem_10_25 (\REG.mem_10_25 ), 
            .n5942(n5942), .\REG.mem_10_24 (\REG.mem_10_24 ), .n5611(n5611), 
            .\REG.mem_6_24 (\REG.mem_6_24 ), .\REG.mem_7_24 (\REG.mem_7_24 ), 
            .\REG.mem_5_24 (\REG.mem_5_24 ), .\REG.mem_4_24 (\REG.mem_4_24 ), 
            .\REG.mem_1_4 (\REG.mem_1_4 ), .\REG.mem_9_24 (\REG.mem_9_24 ), 
            .\REG.mem_8_24 (\REG.mem_8_24 ), .\REG.mem_6_0 (\REG.mem_6_0 ), 
            .\REG.mem_7_0 (\REG.mem_7_0 ), .\REG.mem_5_0 (\REG.mem_5_0 ), 
            .\REG.mem_4_0 (\REG.mem_4_0 ), .\REG.mem_10_4 (\REG.mem_10_4 ), 
            .n5610(n5610), .n5941(n5941), .n5940(n5940), .n5939(n5939), 
            .n5938(n5938), .\REG.mem_10_20 (\REG.mem_10_20 ), .n5937(n5937), 
            .n5608(n5608), .n5604(n5604), .n5603(n5603), .n5602(n5602), 
            .n5936(n5936), .\REG.mem_10_18 (\REG.mem_10_18 ), .n5935(n5935), 
            .n5934(n5934), .\REG.mem_10_16 (\REG.mem_10_16 ), .n5933(n5933), 
            .\REG.mem_1_17 (\REG.mem_1_17 ), .\REG.mem_9_4 (\REG.mem_9_4 ), 
            .\REG.mem_8_4 (\REG.mem_8_4 ), .\REG.mem_6_17 (\REG.mem_6_17 ), 
            .\REG.mem_7_17 (\REG.mem_7_17 ), .\REG.mem_4_17 (\REG.mem_4_17 ), 
            .\REG.mem_5_17 (\REG.mem_5_17 ), .dc32_fifo_read_enable(dc32_fifo_read_enable), 
            .n5932(n5932), .\REG.mem_10_14 (\REG.mem_10_14 ), .n5931(n5931), 
            .n5930(n5930), .\REG.mem_10_12 (\REG.mem_10_12 ), .n5929(n5929), 
            .n5928(n5928), .\REG.mem_10_10 (\REG.mem_10_10 ), .n5927(n5927), 
            .\REG.mem_10_9 (\REG.mem_10_9 ), .n5926(n5926), .n5925(n5925), 
            .\REG.mem_10_7 (\REG.mem_10_7 ), .n5924(n5924), .n5923(n5923), 
            .\REG.mem_10_5 (\REG.mem_10_5 ), .n5922(n5922), .n5921(n5921), 
            .\REG.mem_10_3 (\REG.mem_10_3 ), .n5920(n5920), .n5919(n5919), 
            .\REG.mem_10_1 (\REG.mem_10_1 ), .n5918(n5918), .\REG.mem_10_0 (\REG.mem_10_0 ), 
            .n5917(n5917), .\REG.mem_9_31 (\REG.mem_9_31 ), .n5916(n5916), 
            .\REG.mem_9_30 (\REG.mem_9_30 ), .n5915(n5915), .n5914(n5914), 
            .n5913(n5913), .\REG.mem_9_27 (\REG.mem_9_27 ), .n5912(n5912), 
            .\REG.mem_9_26 (\REG.mem_9_26 ), .n5911(n5911), .\REG.mem_9_25 (\REG.mem_9_25 ), 
            .n5910(n5910), .n5909(n5909), .n5908(n5908), .n5907(n5907), 
            .n5906(n5906), .\REG.mem_9_20 (\REG.mem_9_20 ), .n5905(n5905), 
            .n5904(n5904), .\REG.mem_9_18 (\REG.mem_9_18 ), .n5903(n5903), 
            .n5902(n5902), .\REG.mem_9_16 (\REG.mem_9_16 ), .n5901(n5901), 
            .n5900(n5900), .\REG.mem_9_14 (\REG.mem_9_14 ), .n5899(n5899), 
            .n5898(n5898), .\REG.mem_9_12 (\REG.mem_9_12 ), .n5897(n5897), 
            .n5896(n5896), .\REG.mem_9_10 (\REG.mem_9_10 ), .n5895(n5895), 
            .\REG.mem_9_9 (\REG.mem_9_9 ), .n5894(n5894), .n5893(n5893), 
            .\REG.mem_9_7 (\REG.mem_9_7 ), .n5892(n5892), .n5891(n5891), 
            .n5890(n5890), .n5889(n5889), .\REG.mem_9_3 (\REG.mem_9_3 ), 
            .n5888(n5888), .n5887(n5887), .\REG.mem_9_1 (\REG.mem_9_1 ), 
            .n5886(n5886), .\REG.mem_9_0 (\REG.mem_9_0 ), .n5885(n5885), 
            .\REG.mem_8_31 (\REG.mem_8_31 ), .n5884(n5884), .\REG.mem_8_30 (\REG.mem_8_30 ), 
            .n5883(n5883), .n5882(n5882), .n5881(n5881), .\REG.mem_8_27 (\REG.mem_8_27 ), 
            .n5880(n5880), .\REG.mem_8_26 (\REG.mem_8_26 ), .n5879(n5879), 
            .\REG.mem_8_25 (\REG.mem_8_25 ), .n5878(n5878), .n5877(n5877), 
            .n5876(n5876), .n5875(n5875), .n5874(n5874), .\REG.mem_8_20 (\REG.mem_8_20 ), 
            .n5873(n5873), .n5872(n5872), .\REG.mem_8_18 (\REG.mem_8_18 ), 
            .n5871(n5871), .n5870(n5870), .\REG.mem_8_16 (\REG.mem_8_16 ), 
            .n5869(n5869), .n5868(n5868), .\REG.mem_8_14 (\REG.mem_8_14 ), 
            .n5867(n5867), .n5866(n5866), .\REG.mem_8_12 (\REG.mem_8_12 ), 
            .n5865(n5865), .n5864(n5864), .\REG.mem_8_10 (\REG.mem_8_10 ), 
            .n5863(n5863), .\REG.mem_8_9 (\REG.mem_8_9 ), .n5862(n5862), 
            .n5861(n5861), .\REG.mem_8_7 (\REG.mem_8_7 ), .n5860(n5860), 
            .n5859(n5859), .n5858(n5858), .n5857(n5857), .\REG.mem_8_3 (\REG.mem_8_3 ), 
            .n5856(n5856), .n5855(n5855), .\REG.mem_8_1 (\REG.mem_8_1 ), 
            .n5854(n5854), .\REG.mem_8_0 (\REG.mem_8_0 ), .n5853(n5853), 
            .n5852(n5852), .n5851(n5851), .\REG.mem_7_29 (\REG.mem_7_29 ), 
            .n5850(n5850), .n5849(n5849), .n5848(n5848), .\REG.mem_7_26 (\REG.mem_7_26 ), 
            .n5847(n5847), .\REG.mem_7_25 (\REG.mem_7_25 ), .n5846(n5846), 
            .n5845(n5845), .n5844(n5844), .n5843(n5843), .n5842(n5842), 
            .\REG.mem_7_20 (\REG.mem_7_20 ), .n5841(n5841), .n5840(n5840), 
            .n5839(n5839), .n5838(n5838), .n5837(n5837), .\REG.mem_7_15 (\REG.mem_7_15 ), 
            .n5836(n5836), .\REG.mem_7_14 (\REG.mem_7_14 ), .n5835(n5835), 
            .n5834(n5834), .\REG.mem_7_12 (\REG.mem_7_12 ), .n5833(n5833), 
            .\REG.mem_7_11 (\REG.mem_7_11 ), .n5832(n5832), .n5831(n5831), 
            .n5830(n5830), .\REG.mem_7_8 (\REG.mem_7_8 ), .n5829(n5829), 
            .n5828(n5828), .n5827(n5827), .\REG.mem_7_5 (\REG.mem_7_5 ), 
            .n5826(n5826), .n5825(n5825), .\REG.mem_7_3 (\REG.mem_7_3 ), 
            .n5824(n5824), .n5823(n5823), .n5822(n5822), .n5821(n5821), 
            .n5820(n5820), .n5819(n5819), .\REG.mem_6_29 (\REG.mem_6_29 ), 
            .n5818(n5818), .n5817(n5817), .n5816(n5816), .\REG.mem_6_26 (\REG.mem_6_26 ), 
            .n5815(n5815), .\REG.mem_6_25 (\REG.mem_6_25 ), .n5814(n5814), 
            .n5813(n5813), .n5812(n5812), .n5811(n5811), .n5810(n5810), 
            .\REG.mem_6_20 (\REG.mem_6_20 ), .n5809(n5809), .n5808(n5808), 
            .n5807(n5807), .n5806(n5806), .n5805(n5805), .\REG.mem_6_15 (\REG.mem_6_15 ), 
            .n5804(n5804), .\REG.mem_6_14 (\REG.mem_6_14 ), .n5803(n5803), 
            .n5802(n5802), .\REG.mem_6_12 (\REG.mem_6_12 ), .n5801(n5801), 
            .\REG.mem_6_11 (\REG.mem_6_11 ), .n5800(n5800), .n5799(n5799), 
            .n5798(n5798), .\REG.mem_6_8 (\REG.mem_6_8 ), .n5797(n5797), 
            .n5796(n5796), .n5795(n5795), .\REG.mem_6_5 (\REG.mem_6_5 ), 
            .n5794(n5794), .n5793(n5793), .\REG.mem_6_3 (\REG.mem_6_3 ), 
            .n5792(n5792), .n5791(n5791), .n5790(n5790), .n5789(n5789), 
            .n5788(n5788), .n5600(n5600), .\REG.mem_1_3 (\REG.mem_1_3 ), 
            .n5787(n5787), .\REG.mem_5_29 (\REG.mem_5_29 ), .n25_adj_5(n25_adj_8), 
            .n9(n9), .n5786(n5786), .n5785(n5785), .n5784(n5784), .\REG.mem_5_26 (\REG.mem_5_26 ), 
            .n5783(n5783), .\REG.mem_5_25 (\REG.mem_5_25 ), .n5782(n5782), 
            .\REG.mem_1_16 (\REG.mem_1_16 ), .n5781(n5781), .n5780(n5780), 
            .n5779(n5779), .n5778(n5778), .\REG.mem_5_20 (\REG.mem_5_20 ), 
            .n5777(n5777), .n5776(n5776), .n5775(n5775), .n5774(n5774), 
            .n5773(n5773), .\REG.mem_5_15 (\REG.mem_5_15 ), .n5772(n5772), 
            .\REG.mem_5_14 (\REG.mem_5_14 ), .n5771(n5771), .n5770(n5770), 
            .\REG.mem_5_12 (\REG.mem_5_12 ), .n5769(n5769), .\REG.mem_5_11 (\REG.mem_5_11 ), 
            .\REG.mem_1_25 (\REG.mem_1_25 ), .n5768(n5768), .n5767(n5767), 
            .n5766(n5766), .\REG.mem_5_8 (\REG.mem_5_8 ), .n5765(n5765), 
            .n10(n10), .n26(n26), .n5596(n5596), .n5764(n5764), .n5595(n5595), 
            .\REG.mem_1_5 (\REG.mem_1_5 ), .n5594(n5594), .n5593(n5593), 
            .n5590(n5590), .n5589(n5589), .n5588(n5588), .n5587(n5587), 
            .n5763(n5763), .\REG.mem_5_5 (\REG.mem_5_5 ), .\REG.mem_4_26 (\REG.mem_4_26 ), 
            .n5762(n5762), .n5761(n5761), .\REG.mem_5_3 (\REG.mem_5_3 ), 
            .n5760(n5760), .n5759(n5759), .n5586(n5586), .n5758(n5758), 
            .n5757(n5757), .n5756(n5756), .n5755(n5755), .\REG.mem_4_29 (\REG.mem_4_29 ), 
            .\wr_addr_nxt_c[4] (\wr_addr_nxt_c[4] ), .n5754(n5754), .n5753(n5753), 
            .n5752(n5752), .n5751(n5751), .\REG.mem_4_25 (\REG.mem_4_25 ), 
            .n5750(n5750), .n5749(n5749), .n5748(n5748), .n5747(n5747), 
            .n5585(n5585), .\REG.mem_1_29 (\REG.mem_1_29 ), .n5583(n5583), 
            .n5582(n5582), .n5581(n5581), .\REG.mem_1_8 (\REG.mem_1_8 ), 
            .n5580(n5580), .n5577(n5577), .n5746(n5746), .\REG.mem_4_20 (\REG.mem_4_20 ), 
            .n5745(n5745), .n5744(n5744), .n5743(n5743), .n5742(n5742), 
            .n5741(n5741), .\REG.mem_4_15 (\REG.mem_4_15 ), .n5740(n5740), 
            .\REG.mem_4_14 (\REG.mem_4_14 ), .n5739(n5739), .n5738(n5738), 
            .\REG.mem_4_12 (\REG.mem_4_12 ), .n5574(n5574), .n5572(n5572), 
            .n5571(n5571), .\REG.mem_1_11 (\REG.mem_1_11 ), .n5737(n5737), 
            .\REG.mem_4_11 (\REG.mem_4_11 ), .n5736(n5736), .n5735(n5735), 
            .n5734(n5734), .\REG.mem_4_8 (\REG.mem_4_8 ), .n5733(n5733), 
            .n5732(n5732), .n5731(n5731), .\REG.mem_4_5 (\REG.mem_4_5 ), 
            .n5730(n5730), .n5729(n5729), .\REG.mem_4_3 (\REG.mem_4_3 ), 
            .n5567(n5567), .n5565(n5565), .\REG.mem_1_20 (\REG.mem_1_20 ), 
            .n5564(n5564), .\REG.mem_1_12 (\REG.mem_1_12 ), .n5560(n5560), 
            .n5559(n5559), .\REG.mem_1_14 (\REG.mem_1_14 ), .n5558(n5558), 
            .\REG.mem_1_15 (\REG.mem_1_15 ), .n5557(n5557), .n5556(n5556), 
            .n5555(n5555), .n5554(n5554), .n5551(n5551), .n5550(n5550), 
            .n5728(n5728), .n5727(n5727), .n5726(n5726), .n11(n11), 
            .n27(n27)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_dc_32_lut_gen.v(53[33] 72[34])
    
endmodule
//
// Verilog Description of module fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1
//

module fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1 (dc32_fifo_data_in, 
            \REG.mem_1_9 , GND_net, \REG.mem_6_9 , \REG.mem_7_9 , \REG.mem_4_9 , 
            \REG.mem_5_9 , \REG.mem_24_9 , \REG.mem_25_9 , \REG.mem_1_31 , 
            \REG.mem_9_5 , \REG.mem_8_5 , \REG.mem_26_9 , \REG.mem_27_9 , 
            rd_grey_sync_r, \REG.mem_17_25 , \REG.mem_6_16 , \REG.mem_7_16 , 
            \REG.mem_1_7 , \REG.mem_6_7 , \REG.mem_7_7 , \REG.mem_4_7 , 
            \REG.mem_5_7 , \REG.mem_10_23 , \REG.mem_11_23 , \REG.mem_5_16 , 
            \REG.mem_4_16 , \REG.mem_17_7 , \REG.mem_22_7 , \REG.mem_23_7 , 
            \REG.mem_20_7 , \REG.mem_21_7 , \REG.mem_9_23 , \REG.mem_8_23 , 
            n7, n23, FIFO_CLK_c, DEBUG_1_c, reset_per_frame, wr_fifo_en_w, 
            \wr_addr_r[0] , \REG.mem_22_29 , \REG.mem_23_29 , \REG.mem_21_29 , 
            \REG.mem_20_29 , DEBUG_5_c_0, SLM_CLK_c, \REG.mem_26_21 , 
            \REG.mem_27_21 , \REG.mem_26_25 , \REG.mem_27_25 , \REG.mem_25_25 , 
            \REG.mem_24_25 , \REG.mem_25_21 , \REG.mem_24_21 , \REG.mem_1_10 , 
            \REG.mem_6_10 , \REG.mem_7_10 , \REG.mem_4_10 , \REG.mem_5_10 , 
            \REG.mem_1_26 , n28, n12, dc32_fifo_empty, \wr_grey_sync_r[0] , 
            \aempty_flag_impl.ae_flag_nxt_w , dc32_fifo_almost_empty, n32, 
            n16, \REG.mem_17_10 , \REG.mem_22_10 , \REG.mem_23_10 , 
            \REG.mem_20_10 , \REG.mem_21_10 , dc32_fifo_full, \REG.mem_10_28 , 
            \REG.mem_11_28 , \REG.mem_9_28 , \REG.mem_8_28 , \REG.mem_17_29 , 
            \rd_addr_nxt_c_5__N_573[3] , \rd_addr_nxt_c_5__N_573[1] , n6, 
            n22, \REG.mem_1_28 , \REG.mem_6_28 , \REG.mem_7_28 , \REG.mem_4_28 , 
            \REG.mem_5_28 , \REG.mem_1_2 , \REG.mem_6_2 , \REG.mem_7_2 , 
            \REG.mem_4_2 , \REG.mem_5_2 , \REG.mem_1_22 , \REG.mem_6_22 , 
            \REG.mem_7_22 , \REG.mem_4_22 , \REG.mem_5_22 , \REG.mem_17_22 , 
            \REG.mem_22_22 , \REG.mem_23_22 , \REG.mem_20_22 , \REG.mem_21_22 , 
            \rd_addr_nxt_c_5__N_573[4] , \REG.mem_5_18 , \REG.mem_4_18 , 
            \REG.mem_6_4 , \REG.mem_7_4 , \REG.mem_6_18 , \REG.mem_7_18 , 
            \REG.mem_10_8 , \REG.mem_11_8 , \REG.mem_9_8 , \REG.mem_8_8 , 
            \REG.mem_5_4 , \REG.mem_4_4 , \REG.mem_1_21 , n7013, n7012, 
            n7011, n7010, n7009, n7008, wp_sync1_r, n7007, n7006, 
            n7005, n7004, n7003, n7002, n7000, n6998, n6997, n6996, 
            n6995, n6994, n6993, rp_sync1_r, n6992, n6991, n6990, 
            n6989, \REG.mem_1_13 , n6930, n6928, \wr_addr_r[5] , \REG.mem_6_30 , 
            \REG.mem_7_30 , n6493, \REG.mem_27_31 , n6492, \REG.mem_27_30 , 
            n6491, \REG.mem_27_29 , n6490, \REG.mem_27_28 , n6489, 
            \REG.mem_27_27 , n6488, \REG.mem_27_26 , n6487, n6486, 
            \REG.mem_27_24 , n6485, \REG.mem_27_23 , n6484, \REG.mem_27_22 , 
            n6483, n6482, \REG.mem_27_20 , n6481, \REG.mem_27_19 , 
            n6480, \REG.mem_27_18 , n6479, \REG.mem_27_17 , n6478, 
            \REG.mem_27_16 , n6477, \REG.mem_27_15 , n6476, \REG.mem_27_14 , 
            n6475, \REG.mem_27_13 , n6474, \REG.mem_27_12 , n6473, 
            \REG.mem_27_11 , n6472, \REG.mem_27_10 , n6471, n6470, 
            \REG.mem_27_8 , n6469, \REG.mem_27_7 , n6468, \REG.mem_27_6 , 
            n6467, \REG.mem_27_5 , n6466, \REG.mem_27_4 , n6465, \REG.mem_27_3 , 
            n6464, \REG.mem_27_2 , n6463, \REG.mem_27_1 , n6462, \REG.mem_27_0 , 
            n6461, \REG.mem_26_31 , n6460, \REG.mem_26_30 , n6459, 
            \REG.mem_26_29 , n6458, \REG.mem_26_28 , n6457, \REG.mem_26_27 , 
            n6456, \REG.mem_26_26 , n6455, n6454, \REG.mem_26_24 , 
            n6453, \REG.mem_26_23 , n6452, \REG.mem_26_22 , n6451, 
            n6450, \REG.mem_26_20 , n6449, \REG.mem_26_19 , n6448, 
            \REG.mem_26_18 , n6447, \REG.mem_26_17 , n6446, \REG.mem_26_16 , 
            n6445, \REG.mem_26_15 , n6444, \REG.mem_26_14 , n6443, 
            \REG.mem_26_13 , n6442, \REG.mem_26_12 , n6441, \REG.mem_26_11 , 
            n6440, \REG.mem_26_10 , n6439, n6438, \REG.mem_26_8 , 
            n6437, \REG.mem_26_7 , n6436, \REG.mem_26_6 , n6435, \REG.mem_26_5 , 
            n6434, \REG.mem_26_4 , n6433, \REG.mem_26_3 , n6432, \REG.mem_26_2 , 
            n6431, \REG.mem_26_1 , n6430, \REG.mem_26_0 , n6429, \REG.mem_25_31 , 
            n6428, \REG.mem_25_30 , n6427, \REG.mem_25_29 , n6426, 
            \REG.mem_25_28 , n6425, \REG.mem_25_27 , n6424, \REG.mem_25_26 , 
            n6423, n6422, \REG.mem_25_24 , n6421, \REG.mem_25_23 , 
            n6420, \REG.mem_25_22 , n6419, n6418, \REG.mem_25_20 , 
            n6417, \REG.mem_25_19 , n6416, \REG.mem_25_18 , n6415, 
            \REG.mem_25_17 , n6414, \REG.mem_25_16 , n6413, \REG.mem_25_15 , 
            n6412, \REG.mem_25_14 , n6411, \REG.mem_25_13 , n6410, 
            \REG.mem_25_12 , n6409, \REG.mem_25_11 , n6408, \REG.mem_25_10 , 
            n6407, n6406, \REG.mem_25_8 , n6405, \REG.mem_25_7 , n6404, 
            \REG.mem_25_6 , n6403, \REG.mem_25_5 , n6402, \REG.mem_25_4 , 
            n6401, \REG.mem_25_3 , n6400, \REG.mem_25_2 , n6399, \REG.mem_25_1 , 
            n6398, \REG.mem_25_0 , n6397, \REG.mem_24_31 , n6396, 
            \REG.mem_24_30 , n6395, \REG.mem_24_29 , n6394, \REG.mem_24_28 , 
            n6393, \REG.mem_24_27 , n6392, \REG.mem_24_26 , n6391, 
            n6390, \REG.mem_24_24 , n6389, \REG.mem_24_23 , n6388, 
            \REG.mem_24_22 , n6387, n6386, \REG.mem_24_20 , n6385, 
            \REG.mem_24_19 , n6384, \REG.mem_24_18 , n6383, \REG.mem_24_17 , 
            n6382, \REG.mem_24_16 , n6381, \REG.mem_24_15 , n6380, 
            \REG.mem_24_14 , n6379, \REG.mem_24_13 , n6378, \REG.mem_24_12 , 
            n6377, \REG.mem_24_11 , n6376, \REG.mem_24_10 , n6375, 
            n6374, \REG.mem_24_8 , n6373, \REG.mem_24_7 , n6372, \REG.mem_24_6 , 
            n6371, \REG.mem_24_5 , n6370, \REG.mem_24_4 , n6369, \REG.mem_24_3 , 
            n6368, \REG.mem_24_2 , n6367, \REG.mem_24_1 , n6366, \REG.mem_24_0 , 
            n6365, \REG.mem_23_31 , n6364, \REG.mem_23_30 , n6363, 
            n6362, \REG.mem_23_28 , n6361, \REG.mem_23_27 , n6360, 
            \REG.mem_23_26 , n6359, \REG.mem_23_25 , n6358, \REG.mem_23_24 , 
            n6357, \REG.mem_23_23 , n6356, n6355, \REG.mem_23_21 , 
            n6354, \REG.mem_23_20 , n6353, \REG.mem_23_19 , n6352, 
            \REG.mem_23_18 , n6351, \REG.mem_23_17 , n6350, \REG.mem_23_16 , 
            n6349, \REG.mem_23_15 , n6348, \REG.mem_23_14 , n6347, 
            \REG.mem_23_13 , n6346, \REG.mem_23_12 , n6345, \REG.mem_23_11 , 
            n6344, n6343, \REG.mem_23_9 , n6342, \REG.mem_23_8 , n6341, 
            n6340, \REG.mem_23_6 , n6339, \REG.mem_23_5 , n6338, \REG.mem_23_4 , 
            n6337, \REG.mem_23_3 , n6336, \REG.mem_23_2 , n6335, \REG.mem_23_1 , 
            n6334, \REG.mem_23_0 , n6333, \REG.mem_22_31 , n6332, 
            \REG.mem_22_30 , n6331, n6330, \REG.mem_22_28 , n6329, 
            \REG.mem_22_27 , n6328, \REG.mem_22_26 , n6327, \REG.mem_22_25 , 
            n6326, \REG.mem_22_24 , n6325, \REG.mem_22_23 , n6324, 
            n6323, \REG.mem_22_21 , n6322, \REG.mem_22_20 , n6321, 
            \REG.mem_22_19 , n6320, \REG.mem_22_18 , n6319, \REG.mem_22_17 , 
            n6318, \REG.mem_22_16 , n6317, \REG.mem_22_15 , n6316, 
            \REG.mem_22_14 , n6315, \REG.mem_22_13 , n6314, \REG.mem_22_12 , 
            n6313, \REG.mem_22_11 , n6312, n6311, \REG.mem_22_9 , 
            n6310, \REG.mem_22_8 , n6309, n6308, \REG.mem_22_6 , n6307, 
            \REG.mem_22_5 , n6306, \REG.mem_22_4 , n6305, \REG.mem_22_3 , 
            n6304, \REG.mem_22_2 , n6303, \REG.mem_22_1 , n6302, \REG.mem_22_0 , 
            n6301, \REG.mem_21_31 , n6300, \REG.mem_21_30 , n6299, 
            n6298, \REG.mem_21_28 , n6297, \REG.mem_21_27 , n6296, 
            \REG.mem_21_26 , n6295, \REG.mem_21_25 , n6294, \REG.mem_21_24 , 
            n6293, \REG.mem_21_23 , n6292, n6291, \REG.mem_21_21 , 
            n6290, \REG.mem_21_20 , n6289, \REG.mem_21_19 , n6288, 
            \REG.mem_21_18 , n6287, \REG.mem_21_17 , n6286, \REG.mem_21_16 , 
            n6285, \REG.mem_21_15 , n6284, \REG.mem_21_14 , n6283, 
            \REG.mem_21_13 , n6282, \REG.mem_21_12 , n6281, \REG.mem_21_11 , 
            n6280, n6279, \REG.mem_21_9 , n6278, \REG.mem_21_8 , n6277, 
            n6276, \REG.mem_21_6 , n6275, \REG.mem_21_5 , n6274, \REG.mem_21_4 , 
            n6273, \REG.mem_21_3 , n6272, \REG.mem_21_2 , n6271, \REG.mem_21_1 , 
            n6270, \REG.mem_21_0 , n6269, \REG.mem_20_31 , n6268, 
            \REG.mem_20_30 , n6267, n6266, \REG.mem_20_28 , n6265, 
            \REG.mem_20_27 , n6264, \REG.mem_20_26 , n6263, \REG.mem_20_25 , 
            n6262, \REG.mem_20_24 , n6261, \REG.mem_20_23 , n6260, 
            n6259, \REG.mem_20_21 , n6258, \REG.mem_20_20 , n6257, 
            \REG.mem_20_19 , n6256, \REG.mem_20_18 , n6255, \REG.mem_20_17 , 
            n6254, \REG.mem_20_16 , n6253, \REG.mem_20_15 , n6252, 
            \REG.mem_20_14 , n6251, \REG.mem_20_13 , n6250, \REG.mem_20_12 , 
            n6249, \REG.mem_20_11 , n6248, n6247, \REG.mem_20_9 , 
            n6246, \REG.mem_20_8 , n6245, n6244, \REG.mem_20_6 , n6243, 
            \REG.mem_20_5 , n6242, \REG.mem_20_4 , n6241, \REG.mem_20_3 , 
            n6240, \REG.mem_20_2 , n6239, \REG.mem_20_1 , n6238, \REG.mem_20_0 , 
            n6173, \REG.mem_17_31 , n6172, \REG.mem_17_30 , n6171, 
            n6170, \REG.mem_17_28 , n6169, \REG.mem_17_27 , n6168, 
            \REG.mem_17_26 , n6167, n6166, \REG.mem_17_24 , n6165, 
            \REG.mem_17_23 , n6164, n6163, \REG.mem_17_21 , n6162, 
            \REG.mem_17_20 , n6161, \REG.mem_17_19 , n6160, \REG.mem_17_18 , 
            n6159, \REG.mem_17_17 , n6158, \REG.mem_17_16 , n6157, 
            \REG.mem_17_15 , n6156, \REG.mem_17_14 , n6155, \REG.mem_17_13 , 
            n6154, \REG.mem_17_12 , n6153, \REG.mem_17_11 , n6152, 
            n6151, \REG.mem_17_9 , n6150, \REG.mem_17_8 , n6149, n6148, 
            \REG.mem_17_6 , n6147, \REG.mem_17_5 , n6146, \REG.mem_17_4 , 
            n6145, \REG.mem_17_3 , n6144, \REG.mem_17_2 , n6143, \REG.mem_17_1 , 
            n6142, \REG.mem_17_0 , \REG.mem_5_30 , \REG.mem_4_30 , \REG.mem_1_1 , 
            \REG.mem_6_1 , \REG.mem_7_1 , \REG.mem_4_1 , \REG.mem_5_1 , 
            \REG.mem_6_21 , \REG.mem_7_21 , \REG.mem_5_21 , \REG.mem_4_21 , 
            \REG.mem_1_30 , \REG.mem_10_21 , \REG.mem_11_21 , \REG.mem_1_19 , 
            \REG.mem_6_19 , \REG.mem_7_19 , \REG.mem_5_19 , \REG.mem_4_19 , 
            \REG.mem_9_21 , \REG.mem_8_21 , \wr_addr_p1_w[0] , \REG.mem_6_13 , 
            \REG.mem_7_13 , \REG.mem_5_13 , \REG.mem_4_13 , \REG.mem_10_13 , 
            \REG.mem_11_13 , \REG.mem_9_13 , \REG.mem_8_13 , \REG.mem_10_19 , 
            \REG.mem_11_19 , \REG.mem_9_19 , \REG.mem_8_19 , \REG.mem_1_27 , 
            \REG.mem_6_27 , \REG.mem_7_27 , \REG.mem_4_27 , \REG.mem_5_27 , 
            \REG.mem_1_6 , \REG.mem_8_2 , \REG.mem_9_2 , \REG.mem_10_2 , 
            \REG.mem_11_2 , \wr_addr_nxt_c[2] , VCC_net, dc32_fifo_write_enable, 
            \REG.mem_1_0 , \REG.mem_10_15 , \REG.mem_11_15 , \REG.mem_9_15 , 
            \REG.mem_8_15 , \dc32_fifo_data_out[1] , \REG.mem_10_11 , 
            \REG.mem_11_11 , \REG.mem_9_11 , \REG.mem_8_11 , \dc32_fifo_data_out[2] , 
            \dc32_fifo_data_out[3] , \dc32_fifo_data_out[4] , \dc32_fifo_data_out[5] , 
            \dc32_fifo_data_out[6] , \dc32_fifo_data_out[7] , \dc32_fifo_data_out[8] , 
            \dc32_fifo_data_out[9] , \dc32_fifo_data_out[10] , \dc32_fifo_data_out[11] , 
            \dc32_fifo_data_out[12] , \dc32_fifo_data_out[13] , \dc32_fifo_data_out[14] , 
            \dc32_fifo_data_out[15] , \dc32_fifo_data_out[16] , \dc32_fifo_data_out[17] , 
            \dc32_fifo_data_out[18] , \dc32_fifo_data_out[19] , \dc32_fifo_data_out[20] , 
            \dc32_fifo_data_out[21] , \dc32_fifo_data_out[22] , \dc32_fifo_data_out[23] , 
            \dc32_fifo_data_out[24] , \dc32_fifo_data_out[25] , \dc32_fifo_data_out[26] , 
            \dc32_fifo_data_out[27] , \dc32_fifo_data_out[28] , \dc32_fifo_data_out[29] , 
            \dc32_fifo_data_out[30] , \dc32_fifo_data_out[31] , n7_adj_3, 
            n8, n25, n5981, \REG.mem_11_31 , \REG.mem_1_23 , n5980, 
            \REG.mem_11_30 , \REG.mem_6_6 , \REG.mem_7_6 , \REG.mem_5_6 , 
            \REG.mem_4_6 , n5979, \REG.mem_11_29 , \REG.mem_10_29 , 
            n5978, n5977, \REG.mem_11_27 , n5976, \REG.mem_11_26 , 
            n5975, \REG.mem_11_25 , n5974, \REG.mem_11_24 , \REG.mem_9_29 , 
            \REG.mem_8_29 , n5973, n5972, \REG.mem_11_22 , n29, \REG.mem_8_17 , 
            \REG.mem_9_17 , \REG.mem_10_17 , \REG.mem_11_17 , \REG.mem_1_24 , 
            n5971, n5970, \REG.mem_11_20 , \REG.mem_6_31 , \REG.mem_7_31 , 
            \REG.mem_5_31 , \REG.mem_4_31 , \wr_grey_sync_r[1] , n24, 
            n13, n8_adj_4, \REG.mem_6_23 , \REG.mem_7_23 , \REG.mem_5_23 , 
            \REG.mem_4_23 , \REG.mem_10_6 , \REG.mem_11_6 , n5969, \REG.mem_9_6 , 
            \REG.mem_8_6 , \wr_grey_sync_r[2] , \wr_grey_sync_r[3] , \wr_grey_sync_r[4] , 
            n5968, \REG.mem_11_18 , n5967, n5966, \REG.mem_11_16 , 
            n5965, n5964, \REG.mem_11_14 , n5963, n5962, \REG.mem_11_12 , 
            n5961, n5960, \REG.mem_11_10 , n5959, \REG.mem_11_9 , 
            n5958, n5957, \REG.mem_11_7 , n5956, n5955, \REG.mem_11_5 , 
            n5954, \REG.mem_11_4 , n5953, \REG.mem_11_3 , \REG.mem_10_22 , 
            n5952, n5951, \REG.mem_11_1 , n5950, \REG.mem_11_0 , n5949, 
            \REG.mem_10_31 , n5948, \REG.mem_10_30 , n5947, n5946, 
            n5945, \REG.mem_10_27 , \REG.mem_9_22 , \REG.mem_8_22 , 
            n5944, \REG.mem_10_26 , \REG.mem_1_18 , n5943, \REG.mem_10_25 , 
            n5942, \REG.mem_10_24 , n5611, \REG.mem_6_24 , \REG.mem_7_24 , 
            \REG.mem_5_24 , \REG.mem_4_24 , \REG.mem_1_4 , \REG.mem_9_24 , 
            \REG.mem_8_24 , \REG.mem_6_0 , \REG.mem_7_0 , \REG.mem_5_0 , 
            \REG.mem_4_0 , \REG.mem_10_4 , n5610, n5941, n5940, n5939, 
            n5938, \REG.mem_10_20 , n5937, n5608, n5604, n5603, 
            n5602, n5936, \REG.mem_10_18 , n5935, n5934, \REG.mem_10_16 , 
            n5933, \REG.mem_1_17 , \REG.mem_9_4 , \REG.mem_8_4 , \REG.mem_6_17 , 
            \REG.mem_7_17 , \REG.mem_4_17 , \REG.mem_5_17 , dc32_fifo_read_enable, 
            n5932, \REG.mem_10_14 , n5931, n5930, \REG.mem_10_12 , 
            n5929, n5928, \REG.mem_10_10 , n5927, \REG.mem_10_9 , 
            n5926, n5925, \REG.mem_10_7 , n5924, n5923, \REG.mem_10_5 , 
            n5922, n5921, \REG.mem_10_3 , n5920, n5919, \REG.mem_10_1 , 
            n5918, \REG.mem_10_0 , n5917, \REG.mem_9_31 , n5916, \REG.mem_9_30 , 
            n5915, n5914, n5913, \REG.mem_9_27 , n5912, \REG.mem_9_26 , 
            n5911, \REG.mem_9_25 , n5910, n5909, n5908, n5907, n5906, 
            \REG.mem_9_20 , n5905, n5904, \REG.mem_9_18 , n5903, n5902, 
            \REG.mem_9_16 , n5901, n5900, \REG.mem_9_14 , n5899, n5898, 
            \REG.mem_9_12 , n5897, n5896, \REG.mem_9_10 , n5895, \REG.mem_9_9 , 
            n5894, n5893, \REG.mem_9_7 , n5892, n5891, n5890, n5889, 
            \REG.mem_9_3 , n5888, n5887, \REG.mem_9_1 , n5886, \REG.mem_9_0 , 
            n5885, \REG.mem_8_31 , n5884, \REG.mem_8_30 , n5883, n5882, 
            n5881, \REG.mem_8_27 , n5880, \REG.mem_8_26 , n5879, \REG.mem_8_25 , 
            n5878, n5877, n5876, n5875, n5874, \REG.mem_8_20 , n5873, 
            n5872, \REG.mem_8_18 , n5871, n5870, \REG.mem_8_16 , n5869, 
            n5868, \REG.mem_8_14 , n5867, n5866, \REG.mem_8_12 , n5865, 
            n5864, \REG.mem_8_10 , n5863, \REG.mem_8_9 , n5862, n5861, 
            \REG.mem_8_7 , n5860, n5859, n5858, n5857, \REG.mem_8_3 , 
            n5856, n5855, \REG.mem_8_1 , n5854, \REG.mem_8_0 , n5853, 
            n5852, n5851, \REG.mem_7_29 , n5850, n5849, n5848, \REG.mem_7_26 , 
            n5847, \REG.mem_7_25 , n5846, n5845, n5844, n5843, n5842, 
            \REG.mem_7_20 , n5841, n5840, n5839, n5838, n5837, \REG.mem_7_15 , 
            n5836, \REG.mem_7_14 , n5835, n5834, \REG.mem_7_12 , n5833, 
            \REG.mem_7_11 , n5832, n5831, n5830, \REG.mem_7_8 , n5829, 
            n5828, n5827, \REG.mem_7_5 , n5826, n5825, \REG.mem_7_3 , 
            n5824, n5823, n5822, n5821, n5820, n5819, \REG.mem_6_29 , 
            n5818, n5817, n5816, \REG.mem_6_26 , n5815, \REG.mem_6_25 , 
            n5814, n5813, n5812, n5811, n5810, \REG.mem_6_20 , n5809, 
            n5808, n5807, n5806, n5805, \REG.mem_6_15 , n5804, \REG.mem_6_14 , 
            n5803, n5802, \REG.mem_6_12 , n5801, \REG.mem_6_11 , n5800, 
            n5799, n5798, \REG.mem_6_8 , n5797, n5796, n5795, \REG.mem_6_5 , 
            n5794, n5793, \REG.mem_6_3 , n5792, n5791, n5790, n5789, 
            n5788, n5600, \REG.mem_1_3 , n5787, \REG.mem_5_29 , n25_adj_5, 
            n9, n5786, n5785, n5784, \REG.mem_5_26 , n5783, \REG.mem_5_25 , 
            n5782, \REG.mem_1_16 , n5781, n5780, n5779, n5778, \REG.mem_5_20 , 
            n5777, n5776, n5775, n5774, n5773, \REG.mem_5_15 , n5772, 
            \REG.mem_5_14 , n5771, n5770, \REG.mem_5_12 , n5769, \REG.mem_5_11 , 
            \REG.mem_1_25 , n5768, n5767, n5766, \REG.mem_5_8 , n5765, 
            n10, n26, n5596, n5764, n5595, \REG.mem_1_5 , n5594, 
            n5593, n5590, n5589, n5588, n5587, n5763, \REG.mem_5_5 , 
            \REG.mem_4_26 , n5762, n5761, \REG.mem_5_3 , n5760, n5759, 
            n5586, n5758, n5757, n5756, n5755, \REG.mem_4_29 , \wr_addr_nxt_c[4] , 
            n5754, n5753, n5752, n5751, \REG.mem_4_25 , n5750, n5749, 
            n5748, n5747, n5585, \REG.mem_1_29 , n5583, n5582, n5581, 
            \REG.mem_1_8 , n5580, n5577, n5746, \REG.mem_4_20 , n5745, 
            n5744, n5743, n5742, n5741, \REG.mem_4_15 , n5740, \REG.mem_4_14 , 
            n5739, n5738, \REG.mem_4_12 , n5574, n5572, n5571, \REG.mem_1_11 , 
            n5737, \REG.mem_4_11 , n5736, n5735, n5734, \REG.mem_4_8 , 
            n5733, n5732, n5731, \REG.mem_4_5 , n5730, n5729, \REG.mem_4_3 , 
            n5567, n5565, \REG.mem_1_20 , n5564, \REG.mem_1_12 , n5560, 
            n5559, \REG.mem_1_14 , n5558, \REG.mem_1_15 , n5557, n5556, 
            n5555, n5554, n5551, n5550, n5728, n5727, n5726, n11, 
            n27) /* synthesis syn_module_defined=1 */ ;
    input [31:0]dc32_fifo_data_in;
    output \REG.mem_1_9 ;
    input GND_net;
    output \REG.mem_6_9 ;
    output \REG.mem_7_9 ;
    output \REG.mem_4_9 ;
    output \REG.mem_5_9 ;
    output \REG.mem_24_9 ;
    output \REG.mem_25_9 ;
    output \REG.mem_1_31 ;
    output \REG.mem_9_5 ;
    output \REG.mem_8_5 ;
    output \REG.mem_26_9 ;
    output \REG.mem_27_9 ;
    output [5:0]rd_grey_sync_r;
    output \REG.mem_17_25 ;
    output \REG.mem_6_16 ;
    output \REG.mem_7_16 ;
    output \REG.mem_1_7 ;
    output \REG.mem_6_7 ;
    output \REG.mem_7_7 ;
    output \REG.mem_4_7 ;
    output \REG.mem_5_7 ;
    output \REG.mem_10_23 ;
    output \REG.mem_11_23 ;
    output \REG.mem_5_16 ;
    output \REG.mem_4_16 ;
    output \REG.mem_17_7 ;
    output \REG.mem_22_7 ;
    output \REG.mem_23_7 ;
    output \REG.mem_20_7 ;
    output \REG.mem_21_7 ;
    output \REG.mem_9_23 ;
    output \REG.mem_8_23 ;
    output n7;
    output n23;
    input FIFO_CLK_c;
    output DEBUG_1_c;
    input reset_per_frame;
    output wr_fifo_en_w;
    output \wr_addr_r[0] ;
    output \REG.mem_22_29 ;
    output \REG.mem_23_29 ;
    output \REG.mem_21_29 ;
    output \REG.mem_20_29 ;
    output DEBUG_5_c_0;
    input SLM_CLK_c;
    output \REG.mem_26_21 ;
    output \REG.mem_27_21 ;
    output \REG.mem_26_25 ;
    output \REG.mem_27_25 ;
    output \REG.mem_25_25 ;
    output \REG.mem_24_25 ;
    output \REG.mem_25_21 ;
    output \REG.mem_24_21 ;
    output \REG.mem_1_10 ;
    output \REG.mem_6_10 ;
    output \REG.mem_7_10 ;
    output \REG.mem_4_10 ;
    output \REG.mem_5_10 ;
    output \REG.mem_1_26 ;
    output n28;
    output n12;
    output dc32_fifo_empty;
    output \wr_grey_sync_r[0] ;
    input \aempty_flag_impl.ae_flag_nxt_w ;
    output dc32_fifo_almost_empty;
    output n32;
    output n16;
    output \REG.mem_17_10 ;
    output \REG.mem_22_10 ;
    output \REG.mem_23_10 ;
    output \REG.mem_20_10 ;
    output \REG.mem_21_10 ;
    output dc32_fifo_full;
    output \REG.mem_10_28 ;
    output \REG.mem_11_28 ;
    output \REG.mem_9_28 ;
    output \REG.mem_8_28 ;
    output \REG.mem_17_29 ;
    output \rd_addr_nxt_c_5__N_573[3] ;
    output \rd_addr_nxt_c_5__N_573[1] ;
    output n6;
    output n22;
    output \REG.mem_1_28 ;
    output \REG.mem_6_28 ;
    output \REG.mem_7_28 ;
    output \REG.mem_4_28 ;
    output \REG.mem_5_28 ;
    output \REG.mem_1_2 ;
    output \REG.mem_6_2 ;
    output \REG.mem_7_2 ;
    output \REG.mem_4_2 ;
    output \REG.mem_5_2 ;
    output \REG.mem_1_22 ;
    output \REG.mem_6_22 ;
    output \REG.mem_7_22 ;
    output \REG.mem_4_22 ;
    output \REG.mem_5_22 ;
    output \REG.mem_17_22 ;
    output \REG.mem_22_22 ;
    output \REG.mem_23_22 ;
    output \REG.mem_20_22 ;
    output \REG.mem_21_22 ;
    output \rd_addr_nxt_c_5__N_573[4] ;
    output \REG.mem_5_18 ;
    output \REG.mem_4_18 ;
    output \REG.mem_6_4 ;
    output \REG.mem_7_4 ;
    output \REG.mem_6_18 ;
    output \REG.mem_7_18 ;
    output \REG.mem_10_8 ;
    output \REG.mem_11_8 ;
    output \REG.mem_9_8 ;
    output \REG.mem_8_8 ;
    output \REG.mem_5_4 ;
    output \REG.mem_4_4 ;
    output \REG.mem_1_21 ;
    input n7013;
    input n7012;
    input n7011;
    input n7010;
    input n7009;
    input n7008;
    output [5:0]wp_sync1_r;
    input n7007;
    input n7006;
    input n7005;
    input n7004;
    input n7003;
    input n7002;
    input n7000;
    input n6998;
    input n6997;
    input n6996;
    input n6995;
    input n6994;
    input n6993;
    output [5:0]rp_sync1_r;
    input n6992;
    input n6991;
    input n6990;
    input n6989;
    output \REG.mem_1_13 ;
    input n6930;
    input n6928;
    output \wr_addr_r[5] ;
    output \REG.mem_6_30 ;
    output \REG.mem_7_30 ;
    input n6493;
    output \REG.mem_27_31 ;
    input n6492;
    output \REG.mem_27_30 ;
    input n6491;
    output \REG.mem_27_29 ;
    input n6490;
    output \REG.mem_27_28 ;
    input n6489;
    output \REG.mem_27_27 ;
    input n6488;
    output \REG.mem_27_26 ;
    input n6487;
    input n6486;
    output \REG.mem_27_24 ;
    input n6485;
    output \REG.mem_27_23 ;
    input n6484;
    output \REG.mem_27_22 ;
    input n6483;
    input n6482;
    output \REG.mem_27_20 ;
    input n6481;
    output \REG.mem_27_19 ;
    input n6480;
    output \REG.mem_27_18 ;
    input n6479;
    output \REG.mem_27_17 ;
    input n6478;
    output \REG.mem_27_16 ;
    input n6477;
    output \REG.mem_27_15 ;
    input n6476;
    output \REG.mem_27_14 ;
    input n6475;
    output \REG.mem_27_13 ;
    input n6474;
    output \REG.mem_27_12 ;
    input n6473;
    output \REG.mem_27_11 ;
    input n6472;
    output \REG.mem_27_10 ;
    input n6471;
    input n6470;
    output \REG.mem_27_8 ;
    input n6469;
    output \REG.mem_27_7 ;
    input n6468;
    output \REG.mem_27_6 ;
    input n6467;
    output \REG.mem_27_5 ;
    input n6466;
    output \REG.mem_27_4 ;
    input n6465;
    output \REG.mem_27_3 ;
    input n6464;
    output \REG.mem_27_2 ;
    input n6463;
    output \REG.mem_27_1 ;
    input n6462;
    output \REG.mem_27_0 ;
    input n6461;
    output \REG.mem_26_31 ;
    input n6460;
    output \REG.mem_26_30 ;
    input n6459;
    output \REG.mem_26_29 ;
    input n6458;
    output \REG.mem_26_28 ;
    input n6457;
    output \REG.mem_26_27 ;
    input n6456;
    output \REG.mem_26_26 ;
    input n6455;
    input n6454;
    output \REG.mem_26_24 ;
    input n6453;
    output \REG.mem_26_23 ;
    input n6452;
    output \REG.mem_26_22 ;
    input n6451;
    input n6450;
    output \REG.mem_26_20 ;
    input n6449;
    output \REG.mem_26_19 ;
    input n6448;
    output \REG.mem_26_18 ;
    input n6447;
    output \REG.mem_26_17 ;
    input n6446;
    output \REG.mem_26_16 ;
    input n6445;
    output \REG.mem_26_15 ;
    input n6444;
    output \REG.mem_26_14 ;
    input n6443;
    output \REG.mem_26_13 ;
    input n6442;
    output \REG.mem_26_12 ;
    input n6441;
    output \REG.mem_26_11 ;
    input n6440;
    output \REG.mem_26_10 ;
    input n6439;
    input n6438;
    output \REG.mem_26_8 ;
    input n6437;
    output \REG.mem_26_7 ;
    input n6436;
    output \REG.mem_26_6 ;
    input n6435;
    output \REG.mem_26_5 ;
    input n6434;
    output \REG.mem_26_4 ;
    input n6433;
    output \REG.mem_26_3 ;
    input n6432;
    output \REG.mem_26_2 ;
    input n6431;
    output \REG.mem_26_1 ;
    input n6430;
    output \REG.mem_26_0 ;
    input n6429;
    output \REG.mem_25_31 ;
    input n6428;
    output \REG.mem_25_30 ;
    input n6427;
    output \REG.mem_25_29 ;
    input n6426;
    output \REG.mem_25_28 ;
    input n6425;
    output \REG.mem_25_27 ;
    input n6424;
    output \REG.mem_25_26 ;
    input n6423;
    input n6422;
    output \REG.mem_25_24 ;
    input n6421;
    output \REG.mem_25_23 ;
    input n6420;
    output \REG.mem_25_22 ;
    input n6419;
    input n6418;
    output \REG.mem_25_20 ;
    input n6417;
    output \REG.mem_25_19 ;
    input n6416;
    output \REG.mem_25_18 ;
    input n6415;
    output \REG.mem_25_17 ;
    input n6414;
    output \REG.mem_25_16 ;
    input n6413;
    output \REG.mem_25_15 ;
    input n6412;
    output \REG.mem_25_14 ;
    input n6411;
    output \REG.mem_25_13 ;
    input n6410;
    output \REG.mem_25_12 ;
    input n6409;
    output \REG.mem_25_11 ;
    input n6408;
    output \REG.mem_25_10 ;
    input n6407;
    input n6406;
    output \REG.mem_25_8 ;
    input n6405;
    output \REG.mem_25_7 ;
    input n6404;
    output \REG.mem_25_6 ;
    input n6403;
    output \REG.mem_25_5 ;
    input n6402;
    output \REG.mem_25_4 ;
    input n6401;
    output \REG.mem_25_3 ;
    input n6400;
    output \REG.mem_25_2 ;
    input n6399;
    output \REG.mem_25_1 ;
    input n6398;
    output \REG.mem_25_0 ;
    input n6397;
    output \REG.mem_24_31 ;
    input n6396;
    output \REG.mem_24_30 ;
    input n6395;
    output \REG.mem_24_29 ;
    input n6394;
    output \REG.mem_24_28 ;
    input n6393;
    output \REG.mem_24_27 ;
    input n6392;
    output \REG.mem_24_26 ;
    input n6391;
    input n6390;
    output \REG.mem_24_24 ;
    input n6389;
    output \REG.mem_24_23 ;
    input n6388;
    output \REG.mem_24_22 ;
    input n6387;
    input n6386;
    output \REG.mem_24_20 ;
    input n6385;
    output \REG.mem_24_19 ;
    input n6384;
    output \REG.mem_24_18 ;
    input n6383;
    output \REG.mem_24_17 ;
    input n6382;
    output \REG.mem_24_16 ;
    input n6381;
    output \REG.mem_24_15 ;
    input n6380;
    output \REG.mem_24_14 ;
    input n6379;
    output \REG.mem_24_13 ;
    input n6378;
    output \REG.mem_24_12 ;
    input n6377;
    output \REG.mem_24_11 ;
    input n6376;
    output \REG.mem_24_10 ;
    input n6375;
    input n6374;
    output \REG.mem_24_8 ;
    input n6373;
    output \REG.mem_24_7 ;
    input n6372;
    output \REG.mem_24_6 ;
    input n6371;
    output \REG.mem_24_5 ;
    input n6370;
    output \REG.mem_24_4 ;
    input n6369;
    output \REG.mem_24_3 ;
    input n6368;
    output \REG.mem_24_2 ;
    input n6367;
    output \REG.mem_24_1 ;
    input n6366;
    output \REG.mem_24_0 ;
    input n6365;
    output \REG.mem_23_31 ;
    input n6364;
    output \REG.mem_23_30 ;
    input n6363;
    input n6362;
    output \REG.mem_23_28 ;
    input n6361;
    output \REG.mem_23_27 ;
    input n6360;
    output \REG.mem_23_26 ;
    input n6359;
    output \REG.mem_23_25 ;
    input n6358;
    output \REG.mem_23_24 ;
    input n6357;
    output \REG.mem_23_23 ;
    input n6356;
    input n6355;
    output \REG.mem_23_21 ;
    input n6354;
    output \REG.mem_23_20 ;
    input n6353;
    output \REG.mem_23_19 ;
    input n6352;
    output \REG.mem_23_18 ;
    input n6351;
    output \REG.mem_23_17 ;
    input n6350;
    output \REG.mem_23_16 ;
    input n6349;
    output \REG.mem_23_15 ;
    input n6348;
    output \REG.mem_23_14 ;
    input n6347;
    output \REG.mem_23_13 ;
    input n6346;
    output \REG.mem_23_12 ;
    input n6345;
    output \REG.mem_23_11 ;
    input n6344;
    input n6343;
    output \REG.mem_23_9 ;
    input n6342;
    output \REG.mem_23_8 ;
    input n6341;
    input n6340;
    output \REG.mem_23_6 ;
    input n6339;
    output \REG.mem_23_5 ;
    input n6338;
    output \REG.mem_23_4 ;
    input n6337;
    output \REG.mem_23_3 ;
    input n6336;
    output \REG.mem_23_2 ;
    input n6335;
    output \REG.mem_23_1 ;
    input n6334;
    output \REG.mem_23_0 ;
    input n6333;
    output \REG.mem_22_31 ;
    input n6332;
    output \REG.mem_22_30 ;
    input n6331;
    input n6330;
    output \REG.mem_22_28 ;
    input n6329;
    output \REG.mem_22_27 ;
    input n6328;
    output \REG.mem_22_26 ;
    input n6327;
    output \REG.mem_22_25 ;
    input n6326;
    output \REG.mem_22_24 ;
    input n6325;
    output \REG.mem_22_23 ;
    input n6324;
    input n6323;
    output \REG.mem_22_21 ;
    input n6322;
    output \REG.mem_22_20 ;
    input n6321;
    output \REG.mem_22_19 ;
    input n6320;
    output \REG.mem_22_18 ;
    input n6319;
    output \REG.mem_22_17 ;
    input n6318;
    output \REG.mem_22_16 ;
    input n6317;
    output \REG.mem_22_15 ;
    input n6316;
    output \REG.mem_22_14 ;
    input n6315;
    output \REG.mem_22_13 ;
    input n6314;
    output \REG.mem_22_12 ;
    input n6313;
    output \REG.mem_22_11 ;
    input n6312;
    input n6311;
    output \REG.mem_22_9 ;
    input n6310;
    output \REG.mem_22_8 ;
    input n6309;
    input n6308;
    output \REG.mem_22_6 ;
    input n6307;
    output \REG.mem_22_5 ;
    input n6306;
    output \REG.mem_22_4 ;
    input n6305;
    output \REG.mem_22_3 ;
    input n6304;
    output \REG.mem_22_2 ;
    input n6303;
    output \REG.mem_22_1 ;
    input n6302;
    output \REG.mem_22_0 ;
    input n6301;
    output \REG.mem_21_31 ;
    input n6300;
    output \REG.mem_21_30 ;
    input n6299;
    input n6298;
    output \REG.mem_21_28 ;
    input n6297;
    output \REG.mem_21_27 ;
    input n6296;
    output \REG.mem_21_26 ;
    input n6295;
    output \REG.mem_21_25 ;
    input n6294;
    output \REG.mem_21_24 ;
    input n6293;
    output \REG.mem_21_23 ;
    input n6292;
    input n6291;
    output \REG.mem_21_21 ;
    input n6290;
    output \REG.mem_21_20 ;
    input n6289;
    output \REG.mem_21_19 ;
    input n6288;
    output \REG.mem_21_18 ;
    input n6287;
    output \REG.mem_21_17 ;
    input n6286;
    output \REG.mem_21_16 ;
    input n6285;
    output \REG.mem_21_15 ;
    input n6284;
    output \REG.mem_21_14 ;
    input n6283;
    output \REG.mem_21_13 ;
    input n6282;
    output \REG.mem_21_12 ;
    input n6281;
    output \REG.mem_21_11 ;
    input n6280;
    input n6279;
    output \REG.mem_21_9 ;
    input n6278;
    output \REG.mem_21_8 ;
    input n6277;
    input n6276;
    output \REG.mem_21_6 ;
    input n6275;
    output \REG.mem_21_5 ;
    input n6274;
    output \REG.mem_21_4 ;
    input n6273;
    output \REG.mem_21_3 ;
    input n6272;
    output \REG.mem_21_2 ;
    input n6271;
    output \REG.mem_21_1 ;
    input n6270;
    output \REG.mem_21_0 ;
    input n6269;
    output \REG.mem_20_31 ;
    input n6268;
    output \REG.mem_20_30 ;
    input n6267;
    input n6266;
    output \REG.mem_20_28 ;
    input n6265;
    output \REG.mem_20_27 ;
    input n6264;
    output \REG.mem_20_26 ;
    input n6263;
    output \REG.mem_20_25 ;
    input n6262;
    output \REG.mem_20_24 ;
    input n6261;
    output \REG.mem_20_23 ;
    input n6260;
    input n6259;
    output \REG.mem_20_21 ;
    input n6258;
    output \REG.mem_20_20 ;
    input n6257;
    output \REG.mem_20_19 ;
    input n6256;
    output \REG.mem_20_18 ;
    input n6255;
    output \REG.mem_20_17 ;
    input n6254;
    output \REG.mem_20_16 ;
    input n6253;
    output \REG.mem_20_15 ;
    input n6252;
    output \REG.mem_20_14 ;
    input n6251;
    output \REG.mem_20_13 ;
    input n6250;
    output \REG.mem_20_12 ;
    input n6249;
    output \REG.mem_20_11 ;
    input n6248;
    input n6247;
    output \REG.mem_20_9 ;
    input n6246;
    output \REG.mem_20_8 ;
    input n6245;
    input n6244;
    output \REG.mem_20_6 ;
    input n6243;
    output \REG.mem_20_5 ;
    input n6242;
    output \REG.mem_20_4 ;
    input n6241;
    output \REG.mem_20_3 ;
    input n6240;
    output \REG.mem_20_2 ;
    input n6239;
    output \REG.mem_20_1 ;
    input n6238;
    output \REG.mem_20_0 ;
    input n6173;
    output \REG.mem_17_31 ;
    input n6172;
    output \REG.mem_17_30 ;
    input n6171;
    input n6170;
    output \REG.mem_17_28 ;
    input n6169;
    output \REG.mem_17_27 ;
    input n6168;
    output \REG.mem_17_26 ;
    input n6167;
    input n6166;
    output \REG.mem_17_24 ;
    input n6165;
    output \REG.mem_17_23 ;
    input n6164;
    input n6163;
    output \REG.mem_17_21 ;
    input n6162;
    output \REG.mem_17_20 ;
    input n6161;
    output \REG.mem_17_19 ;
    input n6160;
    output \REG.mem_17_18 ;
    input n6159;
    output \REG.mem_17_17 ;
    input n6158;
    output \REG.mem_17_16 ;
    input n6157;
    output \REG.mem_17_15 ;
    input n6156;
    output \REG.mem_17_14 ;
    input n6155;
    output \REG.mem_17_13 ;
    input n6154;
    output \REG.mem_17_12 ;
    input n6153;
    output \REG.mem_17_11 ;
    input n6152;
    input n6151;
    output \REG.mem_17_9 ;
    input n6150;
    output \REG.mem_17_8 ;
    input n6149;
    input n6148;
    output \REG.mem_17_6 ;
    input n6147;
    output \REG.mem_17_5 ;
    input n6146;
    output \REG.mem_17_4 ;
    input n6145;
    output \REG.mem_17_3 ;
    input n6144;
    output \REG.mem_17_2 ;
    input n6143;
    output \REG.mem_17_1 ;
    input n6142;
    output \REG.mem_17_0 ;
    output \REG.mem_5_30 ;
    output \REG.mem_4_30 ;
    output \REG.mem_1_1 ;
    output \REG.mem_6_1 ;
    output \REG.mem_7_1 ;
    output \REG.mem_4_1 ;
    output \REG.mem_5_1 ;
    output \REG.mem_6_21 ;
    output \REG.mem_7_21 ;
    output \REG.mem_5_21 ;
    output \REG.mem_4_21 ;
    output \REG.mem_1_30 ;
    output \REG.mem_10_21 ;
    output \REG.mem_11_21 ;
    output \REG.mem_1_19 ;
    output \REG.mem_6_19 ;
    output \REG.mem_7_19 ;
    output \REG.mem_5_19 ;
    output \REG.mem_4_19 ;
    output \REG.mem_9_21 ;
    output \REG.mem_8_21 ;
    output \wr_addr_p1_w[0] ;
    output \REG.mem_6_13 ;
    output \REG.mem_7_13 ;
    output \REG.mem_5_13 ;
    output \REG.mem_4_13 ;
    output \REG.mem_10_13 ;
    output \REG.mem_11_13 ;
    output \REG.mem_9_13 ;
    output \REG.mem_8_13 ;
    output \REG.mem_10_19 ;
    output \REG.mem_11_19 ;
    output \REG.mem_9_19 ;
    output \REG.mem_8_19 ;
    output \REG.mem_1_27 ;
    output \REG.mem_6_27 ;
    output \REG.mem_7_27 ;
    output \REG.mem_4_27 ;
    output \REG.mem_5_27 ;
    output \REG.mem_1_6 ;
    output \REG.mem_8_2 ;
    output \REG.mem_9_2 ;
    output \REG.mem_10_2 ;
    output \REG.mem_11_2 ;
    output \wr_addr_nxt_c[2] ;
    input VCC_net;
    input dc32_fifo_write_enable;
    output \REG.mem_1_0 ;
    output \REG.mem_10_15 ;
    output \REG.mem_11_15 ;
    output \REG.mem_9_15 ;
    output \REG.mem_8_15 ;
    output \dc32_fifo_data_out[1] ;
    output \REG.mem_10_11 ;
    output \REG.mem_11_11 ;
    output \REG.mem_9_11 ;
    output \REG.mem_8_11 ;
    output \dc32_fifo_data_out[2] ;
    output \dc32_fifo_data_out[3] ;
    output \dc32_fifo_data_out[4] ;
    output \dc32_fifo_data_out[5] ;
    output \dc32_fifo_data_out[6] ;
    output \dc32_fifo_data_out[7] ;
    output \dc32_fifo_data_out[8] ;
    output \dc32_fifo_data_out[9] ;
    output \dc32_fifo_data_out[10] ;
    output \dc32_fifo_data_out[11] ;
    output \dc32_fifo_data_out[12] ;
    output \dc32_fifo_data_out[13] ;
    output \dc32_fifo_data_out[14] ;
    output \dc32_fifo_data_out[15] ;
    output \dc32_fifo_data_out[16] ;
    output \dc32_fifo_data_out[17] ;
    output \dc32_fifo_data_out[18] ;
    output \dc32_fifo_data_out[19] ;
    output \dc32_fifo_data_out[20] ;
    output \dc32_fifo_data_out[21] ;
    output \dc32_fifo_data_out[22] ;
    output \dc32_fifo_data_out[23] ;
    output \dc32_fifo_data_out[24] ;
    output \dc32_fifo_data_out[25] ;
    output \dc32_fifo_data_out[26] ;
    output \dc32_fifo_data_out[27] ;
    output \dc32_fifo_data_out[28] ;
    output \dc32_fifo_data_out[29] ;
    output \dc32_fifo_data_out[30] ;
    output \dc32_fifo_data_out[31] ;
    output n7_adj_3;
    output n8;
    input n25;
    input n5981;
    output \REG.mem_11_31 ;
    output \REG.mem_1_23 ;
    input n5980;
    output \REG.mem_11_30 ;
    output \REG.mem_6_6 ;
    output \REG.mem_7_6 ;
    output \REG.mem_5_6 ;
    output \REG.mem_4_6 ;
    input n5979;
    output \REG.mem_11_29 ;
    output \REG.mem_10_29 ;
    input n5978;
    input n5977;
    output \REG.mem_11_27 ;
    input n5976;
    output \REG.mem_11_26 ;
    input n5975;
    output \REG.mem_11_25 ;
    input n5974;
    output \REG.mem_11_24 ;
    output \REG.mem_9_29 ;
    output \REG.mem_8_29 ;
    input n5973;
    input n5972;
    output \REG.mem_11_22 ;
    output n29;
    output \REG.mem_8_17 ;
    output \REG.mem_9_17 ;
    output \REG.mem_10_17 ;
    output \REG.mem_11_17 ;
    output \REG.mem_1_24 ;
    input n5971;
    input n5970;
    output \REG.mem_11_20 ;
    output \REG.mem_6_31 ;
    output \REG.mem_7_31 ;
    output \REG.mem_5_31 ;
    output \REG.mem_4_31 ;
    output \wr_grey_sync_r[1] ;
    output n24;
    output n13;
    output n8_adj_4;
    output \REG.mem_6_23 ;
    output \REG.mem_7_23 ;
    output \REG.mem_5_23 ;
    output \REG.mem_4_23 ;
    output \REG.mem_10_6 ;
    output \REG.mem_11_6 ;
    input n5969;
    output \REG.mem_9_6 ;
    output \REG.mem_8_6 ;
    output \wr_grey_sync_r[2] ;
    output \wr_grey_sync_r[3] ;
    output \wr_grey_sync_r[4] ;
    input n5968;
    output \REG.mem_11_18 ;
    input n5967;
    input n5966;
    output \REG.mem_11_16 ;
    input n5965;
    input n5964;
    output \REG.mem_11_14 ;
    input n5963;
    input n5962;
    output \REG.mem_11_12 ;
    input n5961;
    input n5960;
    output \REG.mem_11_10 ;
    input n5959;
    output \REG.mem_11_9 ;
    input n5958;
    input n5957;
    output \REG.mem_11_7 ;
    input n5956;
    input n5955;
    output \REG.mem_11_5 ;
    input n5954;
    output \REG.mem_11_4 ;
    input n5953;
    output \REG.mem_11_3 ;
    output \REG.mem_10_22 ;
    input n5952;
    input n5951;
    output \REG.mem_11_1 ;
    input n5950;
    output \REG.mem_11_0 ;
    input n5949;
    output \REG.mem_10_31 ;
    input n5948;
    output \REG.mem_10_30 ;
    input n5947;
    input n5946;
    input n5945;
    output \REG.mem_10_27 ;
    output \REG.mem_9_22 ;
    output \REG.mem_8_22 ;
    input n5944;
    output \REG.mem_10_26 ;
    output \REG.mem_1_18 ;
    input n5943;
    output \REG.mem_10_25 ;
    input n5942;
    output \REG.mem_10_24 ;
    input n5611;
    output \REG.mem_6_24 ;
    output \REG.mem_7_24 ;
    output \REG.mem_5_24 ;
    output \REG.mem_4_24 ;
    output \REG.mem_1_4 ;
    output \REG.mem_9_24 ;
    output \REG.mem_8_24 ;
    output \REG.mem_6_0 ;
    output \REG.mem_7_0 ;
    output \REG.mem_5_0 ;
    output \REG.mem_4_0 ;
    output \REG.mem_10_4 ;
    input n5610;
    input n5941;
    input n5940;
    input n5939;
    input n5938;
    output \REG.mem_10_20 ;
    input n5937;
    input n5608;
    input n5604;
    input n5603;
    input n5602;
    input n5936;
    output \REG.mem_10_18 ;
    input n5935;
    input n5934;
    output \REG.mem_10_16 ;
    input n5933;
    output \REG.mem_1_17 ;
    output \REG.mem_9_4 ;
    output \REG.mem_8_4 ;
    output \REG.mem_6_17 ;
    output \REG.mem_7_17 ;
    output \REG.mem_4_17 ;
    output \REG.mem_5_17 ;
    input dc32_fifo_read_enable;
    input n5932;
    output \REG.mem_10_14 ;
    input n5931;
    input n5930;
    output \REG.mem_10_12 ;
    input n5929;
    input n5928;
    output \REG.mem_10_10 ;
    input n5927;
    output \REG.mem_10_9 ;
    input n5926;
    input n5925;
    output \REG.mem_10_7 ;
    input n5924;
    input n5923;
    output \REG.mem_10_5 ;
    input n5922;
    input n5921;
    output \REG.mem_10_3 ;
    input n5920;
    input n5919;
    output \REG.mem_10_1 ;
    input n5918;
    output \REG.mem_10_0 ;
    input n5917;
    output \REG.mem_9_31 ;
    input n5916;
    output \REG.mem_9_30 ;
    input n5915;
    input n5914;
    input n5913;
    output \REG.mem_9_27 ;
    input n5912;
    output \REG.mem_9_26 ;
    input n5911;
    output \REG.mem_9_25 ;
    input n5910;
    input n5909;
    input n5908;
    input n5907;
    input n5906;
    output \REG.mem_9_20 ;
    input n5905;
    input n5904;
    output \REG.mem_9_18 ;
    input n5903;
    input n5902;
    output \REG.mem_9_16 ;
    input n5901;
    input n5900;
    output \REG.mem_9_14 ;
    input n5899;
    input n5898;
    output \REG.mem_9_12 ;
    input n5897;
    input n5896;
    output \REG.mem_9_10 ;
    input n5895;
    output \REG.mem_9_9 ;
    input n5894;
    input n5893;
    output \REG.mem_9_7 ;
    input n5892;
    input n5891;
    input n5890;
    input n5889;
    output \REG.mem_9_3 ;
    input n5888;
    input n5887;
    output \REG.mem_9_1 ;
    input n5886;
    output \REG.mem_9_0 ;
    input n5885;
    output \REG.mem_8_31 ;
    input n5884;
    output \REG.mem_8_30 ;
    input n5883;
    input n5882;
    input n5881;
    output \REG.mem_8_27 ;
    input n5880;
    output \REG.mem_8_26 ;
    input n5879;
    output \REG.mem_8_25 ;
    input n5878;
    input n5877;
    input n5876;
    input n5875;
    input n5874;
    output \REG.mem_8_20 ;
    input n5873;
    input n5872;
    output \REG.mem_8_18 ;
    input n5871;
    input n5870;
    output \REG.mem_8_16 ;
    input n5869;
    input n5868;
    output \REG.mem_8_14 ;
    input n5867;
    input n5866;
    output \REG.mem_8_12 ;
    input n5865;
    input n5864;
    output \REG.mem_8_10 ;
    input n5863;
    output \REG.mem_8_9 ;
    input n5862;
    input n5861;
    output \REG.mem_8_7 ;
    input n5860;
    input n5859;
    input n5858;
    input n5857;
    output \REG.mem_8_3 ;
    input n5856;
    input n5855;
    output \REG.mem_8_1 ;
    input n5854;
    output \REG.mem_8_0 ;
    input n5853;
    input n5852;
    input n5851;
    output \REG.mem_7_29 ;
    input n5850;
    input n5849;
    input n5848;
    output \REG.mem_7_26 ;
    input n5847;
    output \REG.mem_7_25 ;
    input n5846;
    input n5845;
    input n5844;
    input n5843;
    input n5842;
    output \REG.mem_7_20 ;
    input n5841;
    input n5840;
    input n5839;
    input n5838;
    input n5837;
    output \REG.mem_7_15 ;
    input n5836;
    output \REG.mem_7_14 ;
    input n5835;
    input n5834;
    output \REG.mem_7_12 ;
    input n5833;
    output \REG.mem_7_11 ;
    input n5832;
    input n5831;
    input n5830;
    output \REG.mem_7_8 ;
    input n5829;
    input n5828;
    input n5827;
    output \REG.mem_7_5 ;
    input n5826;
    input n5825;
    output \REG.mem_7_3 ;
    input n5824;
    input n5823;
    input n5822;
    input n5821;
    input n5820;
    input n5819;
    output \REG.mem_6_29 ;
    input n5818;
    input n5817;
    input n5816;
    output \REG.mem_6_26 ;
    input n5815;
    output \REG.mem_6_25 ;
    input n5814;
    input n5813;
    input n5812;
    input n5811;
    input n5810;
    output \REG.mem_6_20 ;
    input n5809;
    input n5808;
    input n5807;
    input n5806;
    input n5805;
    output \REG.mem_6_15 ;
    input n5804;
    output \REG.mem_6_14 ;
    input n5803;
    input n5802;
    output \REG.mem_6_12 ;
    input n5801;
    output \REG.mem_6_11 ;
    input n5800;
    input n5799;
    input n5798;
    output \REG.mem_6_8 ;
    input n5797;
    input n5796;
    input n5795;
    output \REG.mem_6_5 ;
    input n5794;
    input n5793;
    output \REG.mem_6_3 ;
    input n5792;
    input n5791;
    input n5790;
    input n5789;
    input n5788;
    input n5600;
    output \REG.mem_1_3 ;
    input n5787;
    output \REG.mem_5_29 ;
    output n25_adj_5;
    output n9;
    input n5786;
    input n5785;
    input n5784;
    output \REG.mem_5_26 ;
    input n5783;
    output \REG.mem_5_25 ;
    input n5782;
    output \REG.mem_1_16 ;
    input n5781;
    input n5780;
    input n5779;
    input n5778;
    output \REG.mem_5_20 ;
    input n5777;
    input n5776;
    input n5775;
    input n5774;
    input n5773;
    output \REG.mem_5_15 ;
    input n5772;
    output \REG.mem_5_14 ;
    input n5771;
    input n5770;
    output \REG.mem_5_12 ;
    input n5769;
    output \REG.mem_5_11 ;
    output \REG.mem_1_25 ;
    input n5768;
    input n5767;
    input n5766;
    output \REG.mem_5_8 ;
    input n5765;
    output n10;
    output n26;
    input n5596;
    input n5764;
    input n5595;
    output \REG.mem_1_5 ;
    input n5594;
    input n5593;
    input n5590;
    input n5589;
    input n5588;
    input n5587;
    input n5763;
    output \REG.mem_5_5 ;
    output \REG.mem_4_26 ;
    input n5762;
    input n5761;
    output \REG.mem_5_3 ;
    input n5760;
    input n5759;
    input n5586;
    input n5758;
    input n5757;
    input n5756;
    input n5755;
    output \REG.mem_4_29 ;
    output \wr_addr_nxt_c[4] ;
    input n5754;
    input n5753;
    input n5752;
    input n5751;
    output \REG.mem_4_25 ;
    input n5750;
    input n5749;
    input n5748;
    input n5747;
    input n5585;
    output \REG.mem_1_29 ;
    input n5583;
    input n5582;
    input n5581;
    output \REG.mem_1_8 ;
    input n5580;
    input n5577;
    input n5746;
    output \REG.mem_4_20 ;
    input n5745;
    input n5744;
    input n5743;
    input n5742;
    input n5741;
    output \REG.mem_4_15 ;
    input n5740;
    output \REG.mem_4_14 ;
    input n5739;
    input n5738;
    output \REG.mem_4_12 ;
    input n5574;
    input n5572;
    input n5571;
    output \REG.mem_1_11 ;
    input n5737;
    output \REG.mem_4_11 ;
    input n5736;
    input n5735;
    input n5734;
    output \REG.mem_4_8 ;
    input n5733;
    input n5732;
    input n5731;
    output \REG.mem_4_5 ;
    input n5730;
    input n5729;
    output \REG.mem_4_3 ;
    input n5567;
    input n5565;
    output \REG.mem_1_20 ;
    input n5564;
    output \REG.mem_1_12 ;
    input n5560;
    input n5559;
    output \REG.mem_1_14 ;
    input n5558;
    output \REG.mem_1_15 ;
    input n5557;
    input n5556;
    input n5555;
    input n5554;
    input n5551;
    input n5550;
    input n5728;
    input n5727;
    input n5726;
    output n11;
    output n27;
>>>>>>> Stashed changes
    
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
<<<<<<< Updated upstream
    wire n13875;
    wire [3:0]state_3__N_80;
    
    wire n10833, n10814, n1951;
    wire [31:0]n1880;
    wire [31:0]n1952;
    wire [31:0]n506;
    
    wire n4491;
    wire [31:0]state_timeout_counter;   // src/timing_controller.v(52[12:33])
    
    wire n4809, n12053, n12051, n10121, n10122, n10105, n10106, 
        n12050, n10104, n12043, n10120, n10103, n12044, n10119, 
        n10102, n10118, n12036, n10117, n10132, n10131, n12045, 
        n10116, n12046, n10115, n10130, n10114, n12047, n10113, 
        n10129, n10128, n10127, n10112, n12048, n10111, n10126, 
        n12049, n10110, n10109, n12039, n10125, n12040, n10124, 
        n12041, n10123, n10108;
    wire [3:0]n968;
    
    wire n10107, n4806, n12054, n10823, n12042, n12106, n2033, 
        n4496, n10837, n38, n52, n56, n54, n55, n53, n50, 
        n58, n62, n49, n7570, n7, n12202, n5;
    
    SB_LUT4 i3_4_lut (.I0(state[3]), .I1(state[0]), .I2(state[1]), .I3(state[2]), 
            .O(n13875));
    defparam i3_4_lut.LUT_INIT = 16'h0400;
    SB_DFFE state_i0 (.Q(state[0]), .C(SLM_CLK_c), .E(n10833), .D(state_3__N_80[0]));   // src/timing_controller.v(56[8] 132[4])
    SB_LUT4 mux_898_i25_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[24]), .O(n1952[24]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i25_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i24_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[23]), .O(n1952[23]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i24_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i23_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[22]), .O(n1952[22]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i23_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i21_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[20]), .O(n1952[20]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i21_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i20_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[19]), .O(n1952[19]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i20_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i19_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[18]), .O(n1952[18]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i19_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i16_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[15]), .O(n1952[15]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i16_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i15_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[14]), .O(n1952[14]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i15_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i13_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[12]), .O(n1952[12]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i13_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i10_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[9]), .O(n1952[9]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i10_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i11_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[10]), .O(n1952[10]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i11_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i4_3_lut_4_lut (.I0(state[1]), .I1(n10814), .I2(n1951), 
            .I3(n1880[3]), .O(n1952[3]));   // src/timing_controller.v(56[8] 132[4])
    defparam mux_898_i4_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_DFFESR state_timeout_counter_i0_i31 (.Q(state_timeout_counter[31]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[31]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i30 (.Q(state_timeout_counter[30]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[30]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_LUT4 mux_890_i2_3_lut (.I0(n12053), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[1]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i2_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i3_3_lut (.I0(n12051), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[2]));   // src/timing_controller.v(62[5] 131[12])
    defparam mux_890_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFE state_i3 (.Q(state[3]), .C(SLM_CLK_c), .E(VCC_net), .D(n10514));   // src/timing_controller.v(56[8] 132[4])
    SB_DFF invert_55_i0 (.Q(reset_per_frame), .C(SLM_CLK_c), .D(n10808));   // src/timing_controller.v(62[5] 131[12])
    SB_DFFESR state_timeout_counter_i0_i29 (.Q(state_timeout_counter[29]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[29]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i28 (.Q(state_timeout_counter[28]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[28]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i27 (.Q(state_timeout_counter[27]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[27]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i26 (.Q(state_timeout_counter[26]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[26]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i25 (.Q(state_timeout_counter[25]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[25]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i21 (.Q(state_timeout_counter[21]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[21]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i17 (.Q(state_timeout_counter[17]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[17]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i16 (.Q(state_timeout_counter[16]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[16]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i13 (.Q(state_timeout_counter[13]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[13]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i11 (.Q(state_timeout_counter[11]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[11]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_CARRY sub_31_add_2_22 (.CI(n10121), .I0(state_timeout_counter[20]), 
            .I1(VCC_net), .CO(n10122));
    SB_CARRY sub_31_add_2_6 (.CI(n10105), .I0(state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n10106));
    SB_LUT4 sub_31_add_2_5_lut (.I0(n1774), .I1(state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n10104), .O(n12050)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_21_lut (.I0(n1774), .I1(state_timeout_counter[19]), 
            .I2(VCC_net), .I3(n10120), .O(n12043)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_21 (.CI(n10120), .I0(state_timeout_counter[19]), 
            .I1(VCC_net), .CO(n10121));
    SB_CARRY sub_31_add_2_5 (.CI(n10104), .I0(state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n10105));
    SB_LUT4 sub_31_add_2_4_lut (.I0(n7386), .I1(state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n10103), .O(n12051)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_31_add_2_20_lut (.I0(n1774), .I1(state_timeout_counter[18]), 
            .I2(VCC_net), .I3(n10119), .O(n12044)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_20 (.CI(n10119), .I0(state_timeout_counter[18]), 
            .I1(VCC_net), .CO(n10120));
    SB_CARRY sub_31_add_2_4 (.CI(n10103), .I0(state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n10104));
    SB_LUT4 sub_31_add_2_3_lut (.I0(n1774), .I1(state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n10102), .O(n12053)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_19_lut (.I0(GND_net), .I1(state_timeout_counter[17]), 
            .I2(VCC_net), .I3(n10118), .O(n506[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_19 (.CI(n10118), .I0(state_timeout_counter[17]), 
            .I1(VCC_net), .CO(n10119));
    SB_CARRY sub_31_add_2_3 (.CI(n10102), .I0(state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n10103));
    SB_LUT4 sub_31_add_2_2_lut (.I0(n7386), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n12036)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_31_add_2_18_lut (.I0(GND_net), .I1(state_timeout_counter[16]), 
            .I2(VCC_net), .I3(n10117), .O(n506[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_33_lut (.I0(GND_net), .I1(state_timeout_counter[31]), 
            .I2(VCC_net), .I3(n10132), .O(n506[31])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_32_lut (.I0(GND_net), .I1(state_timeout_counter[30]), 
            .I2(VCC_net), .I3(n10131), .O(n506[30])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_18 (.CI(n10117), .I0(state_timeout_counter[16]), 
            .I1(VCC_net), .CO(n10118));
    SB_CARRY sub_31_add_2_2 (.CI(VCC_net), .I0(state_timeout_counter[0]), 
            .I1(GND_net), .CO(n10102));
    SB_LUT4 sub_31_add_2_17_lut (.I0(n1774), .I1(state_timeout_counter[15]), 
            .I2(VCC_net), .I3(n10116), .O(n12045)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_32 (.CI(n10131), .I0(state_timeout_counter[30]), 
            .I1(VCC_net), .CO(n10132));
    SB_CARRY sub_31_add_2_17 (.CI(n10116), .I0(state_timeout_counter[15]), 
            .I1(VCC_net), .CO(n10117));
    SB_LUT4 sub_31_add_2_16_lut (.I0(n1774), .I1(state_timeout_counter[14]), 
            .I2(VCC_net), .I3(n10115), .O(n12046)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_31_lut (.I0(GND_net), .I1(state_timeout_counter[29]), 
            .I2(VCC_net), .I3(n10130), .O(n506[29])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_16 (.CI(n10115), .I0(state_timeout_counter[14]), 
            .I1(VCC_net), .CO(n10116));
    SB_LUT4 sub_31_add_2_15_lut (.I0(GND_net), .I1(state_timeout_counter[13]), 
            .I2(VCC_net), .I3(n10114), .O(n506[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_31 (.CI(n10130), .I0(state_timeout_counter[29]), 
            .I1(VCC_net), .CO(n10131));
    SB_CARRY sub_31_add_2_15 (.CI(n10114), .I0(state_timeout_counter[13]), 
            .I1(VCC_net), .CO(n10115));
    SB_LUT4 sub_31_add_2_14_lut (.I0(n1774), .I1(state_timeout_counter[12]), 
            .I2(VCC_net), .I3(n10113), .O(n12047)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_30_lut (.I0(GND_net), .I1(state_timeout_counter[28]), 
            .I2(VCC_net), .I3(n10129), .O(n506[28])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_30 (.CI(n10129), .I0(state_timeout_counter[28]), 
            .I1(VCC_net), .CO(n10130));
    SB_LUT4 sub_31_add_2_29_lut (.I0(GND_net), .I1(state_timeout_counter[27]), 
            .I2(VCC_net), .I3(n10128), .O(n506[27])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_29 (.CI(n10128), .I0(state_timeout_counter[27]), 
            .I1(VCC_net), .CO(n10129));
    SB_LUT4 sub_31_add_2_28_lut (.I0(GND_net), .I1(state_timeout_counter[26]), 
            .I2(VCC_net), .I3(n10127), .O(n506[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_14 (.CI(n10113), .I0(state_timeout_counter[12]), 
            .I1(VCC_net), .CO(n10114));
    SB_LUT4 sub_31_add_2_13_lut (.I0(GND_net), .I1(state_timeout_counter[11]), 
            .I2(VCC_net), .I3(n10112), .O(n506[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_28 (.CI(n10127), .I0(state_timeout_counter[26]), 
            .I1(VCC_net), .CO(n10128));
    SB_CARRY sub_31_add_2_13 (.CI(n10112), .I0(state_timeout_counter[11]), 
            .I1(VCC_net), .CO(n10113));
    SB_LUT4 sub_31_add_2_12_lut (.I0(n1774), .I1(state_timeout_counter[10]), 
            .I2(VCC_net), .I3(n10111), .O(n12048)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_27_lut (.I0(GND_net), .I1(state_timeout_counter[25]), 
            .I2(VCC_net), .I3(n10126), .O(n506[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_12 (.CI(n10111), .I0(state_timeout_counter[10]), 
            .I1(VCC_net), .CO(n10112));
    SB_LUT4 sub_31_add_2_11_lut (.I0(n1774), .I1(state_timeout_counter[9]), 
            .I2(VCC_net), .I3(n10110), .O(n12049)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_27 (.CI(n10126), .I0(state_timeout_counter[25]), 
            .I1(VCC_net), .CO(n10127));
    SB_CARRY sub_31_add_2_11 (.CI(n10110), .I0(state_timeout_counter[9]), 
            .I1(VCC_net), .CO(n10111));
    SB_LUT4 sub_31_add_2_10_lut (.I0(GND_net), .I1(state_timeout_counter[8]), 
            .I2(VCC_net), .I3(n10109), .O(n506[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_26_lut (.I0(n1774), .I1(state_timeout_counter[24]), 
            .I2(VCC_net), .I3(n10125), .O(n12039)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_26 (.CI(n10125), .I0(state_timeout_counter[24]), 
            .I1(VCC_net), .CO(n10126));
    SB_LUT4 sub_31_add_2_25_lut (.I0(n1774), .I1(state_timeout_counter[23]), 
            .I2(VCC_net), .I3(n10124), .O(n12040)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_25 (.CI(n10124), .I0(state_timeout_counter[23]), 
            .I1(VCC_net), .CO(n10125));
    SB_LUT4 sub_31_add_2_24_lut (.I0(n1774), .I1(state_timeout_counter[22]), 
            .I2(VCC_net), .I3(n10123), .O(n12041)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_10 (.CI(n10109), .I0(state_timeout_counter[8]), 
            .I1(VCC_net), .CO(n10110));
    SB_LUT4 sub_31_add_2_9_lut (.I0(GND_net), .I1(state_timeout_counter[7]), 
            .I2(VCC_net), .I3(n10108), .O(n506[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_24 (.CI(n10123), .I0(state_timeout_counter[22]), 
            .I1(VCC_net), .CO(n10124));
    SB_DFFESR state_timeout_counter_i0_i8 (.Q(state_timeout_counter[8]), .C(SLM_CLK_c), 
            .E(n4491), .D(n506[8]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFF invert_55_i3 (.Q(INVERT_c_3), .C(SLM_CLK_c), .D(n968[3]));   // src/timing_controller.v(62[5] 131[12])
    SB_CARRY sub_31_add_2_9 (.CI(n10108), .I0(state_timeout_counter[7]), 
            .I1(VCC_net), .CO(n10109));
    SB_LUT4 sub_31_add_2_8_lut (.I0(GND_net), .I1(state_timeout_counter[6]), 
            .I2(VCC_net), .I3(n10107), .O(n506[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_23_lut (.I0(GND_net), .I1(state_timeout_counter[21]), 
            .I2(VCC_net), .I3(n10122), .O(n506[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_8 (.CI(n10107), .I0(state_timeout_counter[6]), 
            .I1(VCC_net), .CO(n10108));
    SB_DFFESR state_timeout_counter_i0_i7 (.Q(state_timeout_counter[7]), .C(SLM_CLK_c), 
            .E(n4491), .D(n506[7]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i6 (.Q(state_timeout_counter[6]), .C(SLM_CLK_c), 
            .E(n4491), .D(n506[6]), .R(n4809));   // src/timing_controller.v(56[8] 132[4])
    SB_DFFESR state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1880[2]), .R(n4806));   // src/timing_controller.v(56[8] 132[4])
>>>>>>> master
    SB_DFFESR state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(SLM_CLK_c), 
            .E(n5068), .D(n630[1]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 i1_2_lut_3_lut (.I0(fifo_state[0]), .I1(DEBUG_8_c), .I2(fifo_state[2]), 
            .I3(GND_net), .O(n7264));   // src/timing_controller.v(88[8] 151[4])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut (.I0(fifo_state[1]), .I1(n11049), .I2(GND_net), .I3(GND_net), 
            .O(n11050));   // src/timing_controller.v(88[8] 151[4])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2620_2_lut (.I0(state[1]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n4070));   // src/timing_controller.v(160[5] 229[12])
    defparam i2620_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_117 (.I0(fifo_state[1]), .I1(fifo_state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6520));   // src/timing_controller.v(88[8] 151[4])
    defparam i1_2_lut_adj_117.LUT_INIT = 16'hdddd;
    SB_LUT4 i12_3_lut_4_lut (.I0(fifo_state[0]), .I1(DEBUG_8_c), .I2(fifo_state[1]), 
            .I3(n40), .O(n3_c));   // src/timing_controller.v(88[8] 151[4])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h8f80;
    SB_LUT4 i1_2_lut_adj_118 (.I0(state[0]), .I1(state[3]), .I2(GND_net), 
            .I3(GND_net), .O(n69));   // src/timing_controller.v(78[11:16])
    defparam i1_2_lut_adj_118.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(fifo_state[2]), .I1(DEBUG_6_c), .I2(n69), .I3(n4070), 
            .O(n4));   // src/timing_controller.v(78[11:16])
    defparam i1_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i5810_4_lut (.I0(n31), .I1(n6520), .I2(fifo_state[0]), .I3(DEBUG_8_c), 
            .O(n7261));   // src/timing_controller.v(77[11:21])
    defparam i5810_4_lut.LUT_INIT = 16'h3505;
    SB_LUT4 sub_71_add_2_26_lut (.I0(GND_net), .I1(state_timeout_counter[24]), 
            .I2(VCC_net), .I3(n10273), .O(n630[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 fifo_state_2__I_0_110_i7_4_lut (.I0(n3_c), .I1(n11406), .I2(fifo_state[2]), 
            .I3(fifo_state[1]), .O(dc32_fifo_read_enable_N_359));   // src/timing_controller.v(93[5] 150[12])
    defparam fifo_state_2__I_0_110_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i5814_3_lut (.I0(n7261), .I1(n7264), .I2(fifo_state[1]), .I3(GND_net), 
            .O(n7265));   // src/timing_controller.v(77[11:21])
    defparam i5814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5818_4_lut (.I0(n4), .I1(n7264), .I2(fifo_state[1]), .I3(fifo_state[0]), 
            .O(n7269));   // src/timing_controller.v(77[11:21])
    defparam i5818_4_lut.LUT_INIT = 16'hcfc5;
    SB_LUT4 i6621_3_lut (.I0(n63), .I1(state[1]), .I2(state[2]), .I3(GND_net), 
            .O(n8067));
    defparam i6621_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_119 (.I0(n5132), .I1(\state_timeout_counter[7] ), 
            .I2(n3), .I3(n11094), .O(n5500));   // src/timing_controller.v(160[5] 229[12])
    defparam i1_4_lut_adj_119.LUT_INIT = 16'ha8a0;
    SB_CARRY sub_71_add_2_26 (.CI(n10273), .I0(state_timeout_counter[24]), 
            .I1(VCC_net), .CO(n10274));
    SB_LUT4 sub_111_add_2_7_lut (.I0(n4_adj_1391), .I1(fifo_state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n10295), .O(n10393)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_120 (.I0(n5132), .I1(n1459), .I2(n106), .I3(n80), 
            .O(n5504));   // src/timing_controller.v(160[5] 229[12])
    defparam i1_4_lut_adj_120.LUT_INIT = 16'ha8a0;
    SB_LUT4 state_3__I_0_105_Mux_0_i7_4_lut (.I0(state[1]), .I1(n63), .I2(state[2]), 
            .I3(state[0]), .O(n7_c));   // src/timing_controller.v(160[5] 229[12])
    defparam state_3__I_0_105_Mux_0_i7_4_lut.LUT_INIT = 16'hc535;
    SB_LUT4 sub_71_add_2_25_lut (.I0(GND_net), .I1(state_timeout_counter[23]), 
            .I2(VCC_net), .I3(n10272), .O(n630[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_3__I_0_105_Mux_0_i15_4_lut (.I0(n7_c), .I1(n8067), .I2(state[3]), 
            .I3(state[0]), .O(state_3__N_83[0]));   // src/timing_controller.v(160[5] 229[12])
    defparam state_3__I_0_105_Mux_0_i15_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 sub_111_add_2_6_lut (.I0(GND_net), .I1(fifo_state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n10294), .O(fifo_state_timeout_counter_5__N_125[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_111_add_2_6 (.CI(n10294), .I0(fifo_state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n10295));
    SB_LUT4 sub_111_add_2_5_lut (.I0(n5), .I1(fifo_state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n10293), .O(n11049)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_5_lut.LUT_INIT = 16'hebbe;
    SB_DFFESR state_timeout_counter_i0_i10 (.Q(state_timeout_counter[10]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[10]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i12 (.Q(state_timeout_counter[12]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[12]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 i3675_1_lut (.I0(buffer_switch_done), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5132));   // src/timing_controller.v(160[5] 229[12])
    defparam i3675_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_111_add_2_5 (.CI(n10293), .I0(fifo_state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n10294));
    SB_LUT4 sub_111_add_2_4_lut (.I0(GND_net), .I1(fifo_state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n10292), .O(fifo_state_timeout_counter_5__N_125[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_111_add_2_4 (.CI(n10292), .I0(fifo_state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n10293));
    SB_CARRY sub_71_add_2_25 (.CI(n10272), .I0(state_timeout_counter[23]), 
            .I1(VCC_net), .CO(n10273));
    SB_CARRY sub_71_add_2_5 (.CI(n10252), .I0(state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n10253));
    SB_LUT4 i1_2_lut_adj_121 (.I0(state[3]), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n11118));
    defparam i1_2_lut_adj_121.LUT_INIT = 16'hbbbb;
    SB_LUT4 sub_71_add_2_24_lut (.I0(GND_net), .I1(state_timeout_counter[22]), 
            .I2(VCC_net), .I3(n10271), .O(n630[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR state_timeout_counter_i0_i23 (.Q(state_timeout_counter[23]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[23]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 i9911_3_lut (.I0(fifo_state[1]), .I1(fifo_state[0]), .I2(fifo_state[2]), 
            .I3(GND_net), .O(fifo_state_2__N_80[1]));   // src/timing_controller.v(93[5] 150[12])
    defparam i9911_3_lut.LUT_INIT = 16'ha6a6;
    SB_LUT4 sub_111_add_2_3_lut (.I0(GND_net), .I1(fifo_state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n10291), .O(fifo_state_timeout_counter_5__N_125[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9921_4_lut (.I0(n11156), .I1(n6461), .I2(fifo_state[2]), 
            .I3(fifo_state[0]), .O(n11352));
    defparam i9921_4_lut.LUT_INIT = 16'h333a;
    SB_LUT4 i49_4_lut (.I0(n11352), .I1(n26), .I2(fifo_state[1]), .I3(fifo_state[2]), 
            .O(n10676));
    defparam i49_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_996_i3_3_lut (.I0(n11379), .I1(state[1]), .I2(n2072), 
            .I3(GND_net), .O(n2073[2]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_996_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFESR state_timeout_counter_i0_i24 (.Q(state_timeout_counter[24]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[24]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 mux_1004_i3_3_lut (.I0(n2073[2]), .I1(n2106), .I2(n2144), 
            .I3(GND_net), .O(n2145[2]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1004_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1004_i4_4_lut (.I0(n11382), .I1(n2106), .I2(n2144), .I3(n2072), 
            .O(n2145[3]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1004_i4_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i9674_4_lut (.I0(n11347), .I1(state[1]), .I2(n2072), .I3(n2144), 
            .O(n2145[4]));   // src/timing_controller.v(160[5] 229[12])
    defparam i9674_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_996_i6_3_lut (.I0(n11378), .I1(state[1]), .I2(n2072), 
            .I3(GND_net), .O(n2073[5]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_996_i6_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFESR state_timeout_counter_i0_i25 (.Q(state_timeout_counter[25]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[25]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 mux_1004_i6_4_lut (.I0(n2073[5]), .I1(n11092), .I2(n2144), 
            .I3(state[1]), .O(n2145[5]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1004_i6_4_lut.LUT_INIT = 16'hfaca;
    SB_CARRY sub_111_add_2_3 (.CI(n10291), .I0(fifo_state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n10292));
    SB_LUT4 mux_996_i7_3_lut (.I0(n11377), .I1(state[1]), .I2(n2072), 
            .I3(GND_net), .O(n2073[6]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_996_i7_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1004_i7_3_lut (.I0(n2073[6]), .I1(n2106), .I2(n2144), 
            .I3(GND_net), .O(n2145[6]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1004_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_996_i8_3_lut (.I0(n11376), .I1(state[1]), .I2(n2072), 
            .I3(GND_net), .O(n2073[7]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_996_i8_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1004_i8_3_lut (.I0(n2073[7]), .I1(n2106), .I2(n2144), 
            .I3(GND_net), .O(n2145[7]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1004_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_996_i9_3_lut (.I0(n11375), .I1(state[1]), .I2(n2072), 
            .I3(GND_net), .O(n2073[8]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_996_i9_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1004_i9_3_lut (.I0(n2073[8]), .I1(n2106), .I2(n2144), 
            .I3(GND_net), .O(n2145[8]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1004_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_111_add_2_2_lut (.I0(GND_net), .I1(fifo_state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(fifo_state_timeout_counter_5__N_125[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_996_i10_3_lut (.I0(n11374), .I1(state[1]), .I2(n2072), 
            .I3(GND_net), .O(n2073[9]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_996_i10_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1004_i10_3_lut (.I0(n2073[9]), .I1(n2106), .I2(n2144), 
            .I3(GND_net), .O(n2145[9]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1004_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_71_add_2_24 (.CI(n10271), .I0(state_timeout_counter[22]), 
            .I1(VCC_net), .CO(n10272));
    SB_LUT4 mux_996_i12_3_lut (.I0(n11373), .I1(state[1]), .I2(n2072), 
            .I3(GND_net), .O(n2073[11]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_996_i12_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1004_i12_3_lut (.I0(n2073[11]), .I1(n2106), .I2(n2144), 
            .I3(GND_net), .O(n2145[11]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1004_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9971_2_lut (.I0(state[2]), .I1(state[3]), .I2(GND_net), .I3(GND_net), 
            .O(n4068));   // src/timing_controller.v(160[5] 229[12])
    defparam i9971_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 sub_71_add_2_23_lut (.I0(GND_net), .I1(state_timeout_counter[21]), 
            .I2(VCC_net), .I3(n10270), .O(n630[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9615_3_lut (.I0(state[1]), .I1(state[3]), .I2(state[0]), 
            .I3(GND_net), .O(n11191));
    defparam i9615_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY sub_71_add_2_23 (.CI(n10270), .I0(state_timeout_counter[21]), 
            .I1(VCC_net), .CO(n10271));
    SB_LUT4 sub_71_add_2_4_lut (.I0(n7836), .I1(state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n10251), .O(n11379)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_4_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_111_add_2_2 (.CI(VCC_net), .I0(fifo_state_timeout_counter[0]), 
            .I1(GND_net), .CO(n10291));
    SB_LUT4 sub_71_add_2_22_lut (.I0(GND_net), .I1(state_timeout_counter[20]), 
            .I2(VCC_net), .I3(n10269), .O(n630[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_22 (.CI(n10269), .I0(state_timeout_counter[20]), 
            .I1(VCC_net), .CO(n10270));
    SB_CARRY sub_71_add_2_4 (.CI(n10251), .I0(state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n10252));
    SB_LUT4 sub_71_add_2_21_lut (.I0(GND_net), .I1(state_timeout_counter[19]), 
            .I2(VCC_net), .I3(n10268), .O(n630[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_21 (.CI(n10268), .I0(state_timeout_counter[19]), 
            .I1(VCC_net), .CO(n10269));
    SB_LUT4 sub_71_add_2_20_lut (.I0(GND_net), .I1(state_timeout_counter[18]), 
            .I2(VCC_net), .I3(n10267), .O(n630[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR state_timeout_counter_i0_i13 (.Q(state_timeout_counter[13]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[13]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i14 (.Q(state_timeout_counter[14]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[14]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_CARRY sub_71_add_2_20 (.CI(n10267), .I0(state_timeout_counter[18]), 
            .I1(VCC_net), .CO(n10268));
    SB_LUT4 sub_71_add_2_19_lut (.I0(GND_net), .I1(state_timeout_counter[17]), 
            .I2(VCC_net), .I3(n10266), .O(n630[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_71_add_2_3_lut (.I0(GND_net), .I1(state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n10250), .O(n630[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF invert_100_i4 (.Q(INVERT_c_4), .C(SLM_CLK_c), .D(n1103[4]));   // src/timing_controller.v(160[5] 229[12])
    SB_LUT4 i1_2_lut_adj_122 (.I0(n63), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_1392));
    defparam i1_2_lut_adj_122.LUT_INIT = 16'heeee;
    SB_CARRY sub_71_add_2_3 (.CI(n10250), .I0(state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n10251));
    SB_LUT4 sub_71_add_2_2_lut (.I0(n7836), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n11358)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_71_add_2_2 (.CI(VCC_net), .I0(state_timeout_counter[0]), 
            .I1(GND_net), .CO(n10250));
    SB_CARRY sub_71_add_2_19 (.CI(n10266), .I0(state_timeout_counter[17]), 
            .I1(VCC_net), .CO(n10267));
    SB_LUT4 sub_71_add_2_18_lut (.I0(GND_net), .I1(state_timeout_counter[16]), 
            .I2(VCC_net), .I3(n10265), .O(n630[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_18 (.CI(n10265), .I0(state_timeout_counter[16]), 
            .I1(VCC_net), .CO(n10266));
    SB_LUT4 state_3__I_0_105_Mux_1_i15_4_lut (.I0(state[0]), .I1(n4_adj_1392), 
            .I2(state[3]), .I3(state[1]), .O(state_3__N_83[1]));   // src/timing_controller.v(160[5] 229[12])
    defparam state_3__I_0_105_Mux_1_i15_4_lut.LUT_INIT = 16'hf51a;
    SB_LUT4 i1_4_lut_adj_123 (.I0(state[1]), .I1(n11118), .I2(state[0]), 
            .I3(state[2]), .O(n5304));
    defparam i1_4_lut_adj_123.LUT_INIT = 16'hcccd;
    SB_LUT4 sub_71_add_2_17_lut (.I0(GND_net), .I1(state_timeout_counter[15]), 
            .I2(VCC_net), .I3(n10264), .O(n630[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_17 (.CI(n10264), .I0(state_timeout_counter[15]), 
            .I1(VCC_net), .CO(n10265));
    SB_LUT4 state_3__I_0_105_Mux_2_i15_4_lut (.I0(state[1]), .I1(state[2]), 
            .I2(state[3]), .I3(state[0]), .O(state_3__N_83[2]));   // src/timing_controller.v(160[5] 229[12])
    defparam state_3__I_0_105_Mux_2_i15_4_lut.LUT_INIT = 16'hc2ce;
    SB_LUT4 i9679_4_lut (.I0(state[2]), .I1(n63), .I2(n11191), .I3(n5068), 
            .O(n11257));
    defparam i9679_4_lut.LUT_INIT = 16'hc8fa;
    SB_LUT4 sub_71_add_2_16_lut (.I0(GND_net), .I1(state_timeout_counter[14]), 
            .I2(VCC_net), .I3(n10263), .O(n630[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_16 (.CI(n10263), .I0(state_timeout_counter[14]), 
            .I1(VCC_net), .CO(n10264));
    SB_LUT4 sub_71_add_2_15_lut (.I0(GND_net), .I1(state_timeout_counter[13]), 
            .I2(VCC_net), .I3(n10262), .O(n630[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51_3_lut (.I0(dc32_fifo_full), .I1(DEBUG_8_c), .I2(fifo_state[0]), 
            .I3(GND_net), .O(n26));
    defparam i51_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_124 (.I0(state[0]), .I1(state[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11101));
    defparam i1_2_lut_adj_124.LUT_INIT = 16'h2222;
    SB_CARRY sub_71_add_2_15 (.CI(n10262), .I0(state_timeout_counter[13]), 
            .I1(VCC_net), .CO(n10263));
    SB_LUT4 i9843_2_lut_3_lut (.I0(state[0]), .I1(n63), .I2(state[1]), 
            .I3(GND_net), .O(n11356));   // src/timing_controller.v(154[8] 230[4])
    defparam i9843_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i9953_3_lut (.I0(n7), .I1(n59), .I2(n6), .I3(GND_net), .O(\aempty_flag_impl.ae_flag_nxt_w ));
    defparam i9953_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 sub_71_add_2_14_lut (.I0(GND_net), .I1(state_timeout_counter[12]), 
            .I2(VCC_net), .I3(n10261), .O(n630[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_14 (.CI(n10261), .I0(state_timeout_counter[12]), 
            .I1(VCC_net), .CO(n10262));
    SB_LUT4 sub_71_add_2_13_lut (.I0(n1967), .I1(state_timeout_counter[11]), 
            .I2(VCC_net), .I3(n10260), .O(n11373)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_71_add_2_13 (.CI(n10260), .I0(state_timeout_counter[11]), 
            .I1(VCC_net), .CO(n10261));
    SB_LUT4 sub_71_add_2_12_lut (.I0(GND_net), .I1(state_timeout_counter[10]), 
            .I2(VCC_net), .I3(n10259), .O(n630[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_12 (.CI(n10259), .I0(state_timeout_counter[10]), 
            .I1(VCC_net), .CO(n10260));
    SB_DFFESR state_timeout_counter_i0_i15 (.Q(state_timeout_counter[15]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[15]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i16 (.Q(state_timeout_counter[16]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[16]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i17 (.Q(state_timeout_counter[17]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[17]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 i6_2_lut (.I0(state_timeout_counter[19]), .I1(state_timeout_counter[21]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // src/timing_controller.v(154[8] 230[4])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut (.I0(state_timeout_counter[22]), .I1(state_timeout_counter[26]), 
            .I2(state_timeout_counter[25]), .I3(state_timeout_counter[28]), 
            .O(n52));   // src/timing_controller.v(154[8] 230[4])
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR state_timeout_counter_i0_i18 (.Q(state_timeout_counter[18]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[18]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 i2_3_lut_4_lut (.I0(fifo_state[0]), .I1(fifo_state[1]), .I2(fifo_state[2]), 
            .I3(DEBUG_8_c), .O(n5496));   // src/timing_controller.v(77[11:21])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i9580_3_lut (.I0(state[3]), .I1(DEBUG_6_c), .I2(n4943), .I3(GND_net), 
            .O(n11156));
    defparam i9580_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 i24_4_lut (.I0(state_timeout_counter[4]), .I1(state_timeout_counter[16]), 
            .I2(state_timeout_counter[8]), .I3(state_timeout_counter[0]), 
            .O(n56));   // src/timing_controller.v(154[8] 230[4])
    defparam i24_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i22_4_lut (.I0(state_timeout_counter[10]), .I1(state_timeout_counter[17]), 
            .I2(state_timeout_counter[12]), .I3(state_timeout_counter[18]), 
            .O(n54));   // src/timing_controller.v(154[8] 230[4])
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(state_timeout_counter[20]), .I1(state_timeout_counter[1]), 
            .I2(state_timeout_counter[24]), .I3(state_timeout_counter[2]), 
            .O(n55));   // src/timing_controller.v(154[8] 230[4])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF invert_100_i2 (.Q(buffer_switch_done), .C(SLM_CLK_c), .D(n11102));   // src/timing_controller.v(160[5] 229[12])
    SB_DFFESR state_timeout_counter_i0_i19 (.Q(state_timeout_counter[19]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[19]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 i47_1_lut (.I0(dc32_fifo_read_enable), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // src/top.v(482[26:47])
    defparam i47_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR state_timeout_counter_i0_i20 (.Q(state_timeout_counter[20]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[20]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 i12_3_lut_3_lut (.I0(fifo_state[0]), .I1(fifo_state[1]), .I2(fifo_state[2]), 
            .I3(GND_net), .O(fifo_state_2__N_80[2]));   // src/timing_controller.v(77[11:21])
    defparam i12_3_lut_3_lut.LUT_INIT = 16'h5858;
    SB_LUT4 i50_3_lut (.I0(n11156), .I1(n6461), .I2(fifo_state[0]), .I3(GND_net), 
            .O(n28));
    defparam i50_3_lut.LUT_INIT = 16'hc5c5;
    SB_DFFE state_i2 (.Q(state[2]), .C(SLM_CLK_c), .E(n5304), .D(state_3__N_83[2]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_i1 (.Q(state[1]), .C(SLM_CLK_c), .E(n5304), .D(state_3__N_83[1]));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 i9994_4_lut (.I0(fifo_state[2]), .I1(n28), .I2(n26), .I3(fifo_state[1]), 
            .O(n23));
    defparam i9994_4_lut.LUT_INIT = 16'hfabb;
    SB_DFFE state_timeout_counter_i0_i11 (.Q(state_timeout_counter[11]), .C(SLM_CLK_c), 
            .E(n5068), .D(n2145[11]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i9 (.Q(state_timeout_counter[9]), .C(SLM_CLK_c), 
            .E(n5068), .D(n2145[9]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i8 (.Q(state_timeout_counter[8]), .C(SLM_CLK_c), 
            .E(n5068), .D(n2145[8]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i7 (.Q(state_timeout_counter[7]), .C(SLM_CLK_c), 
            .E(n5068), .D(n2145[7]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i6 (.Q(state_timeout_counter[6]), .C(SLM_CLK_c), 
            .E(n5068), .D(n2145[6]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i5 (.Q(state_timeout_counter[5]), .C(SLM_CLK_c), 
            .E(n5068), .D(n2145[5]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(SLM_CLK_c), 
            .E(n5068), .D(n2145[4]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(SLM_CLK_c), 
            .E(n5068), .D(n2145[3]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(SLM_CLK_c), 
            .E(n5068), .D(n2145[2]));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFE fifo_state_i2 (.Q(fifo_state[2]), .C(SLM_CLK_c), .E(n10676), 
            .D(fifo_state_2__N_80[2]));   // src/timing_controller.v(88[8] 151[4])
    SB_LUT4 sub_71_add_2_11_lut (.I0(n1967), .I1(state_timeout_counter[9]), 
            .I2(VCC_net), .I3(n10258), .O(n11374)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_11_lut.LUT_INIT = 16'h8228;
    SB_DFFE fifo_state_i1 (.Q(fifo_state[1]), .C(SLM_CLK_c), .E(n23), 
            .D(fifo_state_2__N_80[1]));   // src/timing_controller.v(88[8] 151[4])
    SB_DFFESR state_timeout_counter_i0_i26 (.Q(state_timeout_counter[26]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[26]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 i12_4_lut (.I0(fifo_state[0]), .I1(fifo_state[1]), .I2(fifo_state[2]), 
            .I3(n6461), .O(fifo_state_2__N_80[0]));   // src/timing_controller.v(77[11:21])
    defparam i12_4_lut.LUT_INIT = 16'ha595;
    SB_DFFESR state_timeout_counter_i0_i27 (.Q(state_timeout_counter[27]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[27]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 i4_4_lut (.I0(fifo_state_timeout_counter[3]), .I1(fifo_state_timeout_counter[2]), 
            .I2(fifo_state_timeout_counter[1]), .I3(fifo_state_timeout_counter[5]), 
            .O(n10));   // src/timing_controller.v(88[8] 151[4])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR state_timeout_counter_i0_i28 (.Q(state_timeout_counter[28]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[28]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_LUT4 i5_3_lut (.I0(fifo_state_timeout_counter[0]), .I1(n10), .I2(fifo_state_timeout_counter[4]), 
            .I3(GND_net), .O(n6461));   // src/timing_controller.v(88[8] 151[4])
    defparam i5_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i21_4_lut (.I0(state_timeout_counter[3]), .I1(state_timeout_counter[6]), 
            .I2(state_timeout_counter[5]), .I3(state_timeout_counter[9]), 
            .O(n53));   // src/timing_controller.v(154[8] 230[4])
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR state_timeout_counter_i0_i29 (.Q(state_timeout_counter[29]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[29]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i30 (.Q(state_timeout_counter[30]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[30]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR state_timeout_counter_i0_i31 (.Q(state_timeout_counter[31]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[31]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_DFFESR fifo_state_timeout_counter_i0_i1 (.Q(fifo_state_timeout_counter[1]), 
            .C(SLM_CLK_c), .E(n7269), .D(fifo_state_timeout_counter_5__N_125[1]), 
            .R(n7265));   // src/timing_controller.v(88[8] 151[4])
    SB_DFFESR fifo_state_timeout_counter_i0_i2 (.Q(fifo_state_timeout_counter[2]), 
            .C(SLM_CLK_c), .E(n7269), .D(fifo_state_timeout_counter_5__N_125[2]), 
            .R(n7265));   // src/timing_controller.v(88[8] 151[4])
    SB_DFFESR fifo_state_timeout_counter_i0_i3 (.Q(fifo_state_timeout_counter[3]), 
            .C(SLM_CLK_c), .E(n7269), .D(n11050), .R(n5496));   // src/timing_controller.v(88[8] 151[4])
    SB_DFFESR fifo_state_timeout_counter_i0_i4 (.Q(fifo_state_timeout_counter[4]), 
            .C(SLM_CLK_c), .E(n7269), .D(fifo_state_timeout_counter_5__N_125[4]), 
            .R(n7265));   // src/timing_controller.v(88[8] 151[4])
    SB_DFFESS fifo_state_timeout_counter_i0_i5 (.Q(fifo_state_timeout_counter[5]), 
            .C(SLM_CLK_c), .E(n7269), .D(n10393), .S(n5496));   // src/timing_controller.v(88[8] 151[4])
    SB_LUT4 i18_4_lut (.I0(state_timeout_counter[29]), .I1(state_timeout_counter[7]), 
            .I2(state_timeout_counter[30]), .I3(state_timeout_counter[11]), 
            .O(n50));   // src/timing_controller.v(154[8] 230[4])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY sub_71_add_2_11 (.CI(n10258), .I0(state_timeout_counter[9]), 
            .I1(VCC_net), .CO(n10259));
    SB_LUT4 sub_71_add_2_10_lut (.I0(n1967), .I1(state_timeout_counter[8]), 
            .I2(VCC_net), .I3(n10257), .O(n11375)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i26_4_lut (.I0(state_timeout_counter[13]), .I1(n52), .I2(n38), 
            .I3(state_timeout_counter[14]), .O(n58));   // src/timing_controller.v(154[8] 230[4])
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30_4_lut (.I0(n53), .I1(n55), .I2(n54), .I3(n56), .O(n62));   // src/timing_controller.v(154[8] 230[4])
    defparam i30_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(state_timeout_counter[31]), .I1(state_timeout_counter[23]), 
            .I2(state_timeout_counter[15]), .I3(state_timeout_counter[27]), 
            .O(n49));   // src/timing_controller.v(154[8] 230[4])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31_4_lut (.I0(n49), .I1(n62), .I2(n58), .I3(n50), .O(n63));   // src/timing_controller.v(154[8] 230[4])
    defparam i31_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_71_add_2_33_lut (.I0(GND_net), .I1(state_timeout_counter[31]), 
            .I2(VCC_net), .I3(n10280), .O(n630[31])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_71_add_2_32_lut (.I0(GND_net), .I1(state_timeout_counter[30]), 
            .I2(VCC_net), .I3(n10279), .O(n630[30])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9959_4_lut (.I0(n5068), .I1(n2072), .I2(n1967), .I3(n2144), 
            .O(n5537));
    defparam i9959_4_lut.LUT_INIT = 16'haa8a;
    SB_CARRY sub_71_add_2_32 (.CI(n10279), .I0(state_timeout_counter[30]), 
            .I1(VCC_net), .CO(n10280));
    SB_LUT4 sub_71_add_2_31_lut (.I0(GND_net), .I1(state_timeout_counter[29]), 
            .I2(VCC_net), .I3(n10278), .O(n630[29])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_31_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR state_timeout_counter_i0_i21 (.Q(state_timeout_counter[21]), 
            .C(SLM_CLK_c), .E(n5068), .D(n630[21]), .R(n5537));   // src/timing_controller.v(154[8] 230[4])
    SB_CARRY sub_71_add_2_31 (.CI(n10278), .I0(state_timeout_counter[29]), 
            .I1(VCC_net), .CO(n10279));
    SB_LUT4 i9926_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n11506));   // src/timing_controller.v(160[5] 229[12])
    defparam i9926_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY sub_71_add_2_10 (.CI(n10257), .I0(state_timeout_counter[8]), 
            .I1(VCC_net), .CO(n10258));
    SB_LUT4 i6501_2_lut (.I0(dc32_fifo_full), .I1(fifo_state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // src/timing_controller.v(93[5] 150[12])
    defparam i6501_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 sub_71_add_2_30_lut (.I0(GND_net), .I1(state_timeout_counter[28]), 
            .I2(VCC_net), .I3(n10277), .O(n630[28])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_30 (.CI(n10277), .I0(state_timeout_counter[28]), 
            .I1(VCC_net), .CO(n10278));
    SB_LUT4 sub_71_add_2_9_lut (.I0(n1967), .I1(state_timeout_counter[7]), 
            .I2(VCC_net), .I3(n10256), .O(n11376)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_71_add_2_29_lut (.I0(GND_net), .I1(state_timeout_counter[27]), 
            .I2(VCC_net), .I3(n10276), .O(n630[27])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_29_lut.LUT_INIT = 16'hC33C;
    SB_DFF invert_100_i0 (.Q(reset_all), .C(SLM_CLK_c), .D(n11104));   // src/timing_controller.v(160[5] 229[12])
    SB_CARRY sub_71_add_2_29 (.CI(n10276), .I0(state_timeout_counter[27]), 
            .I1(VCC_net), .CO(n10277));
    SB_LUT4 i1_2_lut_3_lut_adj_125 (.I0(fifo_state[2]), .I1(n6461), .I2(n4), 
            .I3(GND_net), .O(n31));   // src/timing_controller.v(88[8] 151[4])
    defparam i1_2_lut_3_lut_adj_125.LUT_INIT = 16'hf8f8;
    SB_CARRY sub_71_add_2_9 (.CI(n10256), .I0(state_timeout_counter[7]), 
            .I1(VCC_net), .CO(n10257));
    SB_LUT4 sub_71_add_2_8_lut (.I0(n1967), .I1(state_timeout_counter[6]), 
            .I2(VCC_net), .I3(n10255), .O(n11377)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_71_add_2_28_lut (.I0(GND_net), .I1(state_timeout_counter[26]), 
            .I2(VCC_net), .I3(n10275), .O(n630[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_8 (.CI(n10255), .I0(state_timeout_counter[6]), 
            .I1(VCC_net), .CO(n10256));
    SB_LUT4 sub_71_add_2_7_lut (.I0(n1967), .I1(state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n10254), .O(n11378)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_71_add_2_28 (.CI(n10275), .I0(state_timeout_counter[26]), 
            .I1(VCC_net), .CO(n10276));
    SB_LUT4 i9881_2_lut (.I0(fifo_state[0]), .I1(n6461), .I2(GND_net), 
            .I3(GND_net), .O(n11391));
    defparam i9881_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i51_4_lut (.I0(n11391), .I1(n7264), .I2(fifo_state[1]), .I3(fifo_state[2]), 
            .O(sc32_fifo_read_enable_N_366));
    defparam i51_4_lut.LUT_INIT = 16'hcac0;
    SB_CARRY sub_71_add_2_7 (.CI(n10254), .I0(state_timeout_counter[5]), 
            .I1(VCC_net), .CO(n10255));
    SB_DFF invert_100_i1 (.Q(reset_per_frame), .C(SLM_CLK_c), .D(n11700));   // src/timing_controller.v(160[5] 229[12])
    SB_LUT4 sub_71_add_2_6_lut (.I0(n1967), .I1(state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n10253), .O(n11347)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_6_lut.LUT_INIT = 16'h8228;
    SB_DFFESR fifo_state_timeout_counter_i0_i0 (.Q(fifo_state_timeout_counter[0]), 
            .C(SLM_CLK_c), .E(n7269), .D(fifo_state_timeout_counter_5__N_125[0]), 
            .R(n7265));   // src/timing_controller.v(88[8] 151[4])
    SB_LUT4 i6613_2_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(state[2]), 
            .I3(GND_net), .O(n4943));
    defparam i6613_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_126 (.I0(state[0]), .I1(state[3]), .I2(state[1]), 
            .I3(state[2]), .O(n11102));
    defparam i2_3_lut_4_lut_adj_126.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(state[0]), .I1(n63), .I2(state[2]), 
            .I3(state[3]), .O(n11092));   // src/timing_controller.v(154[8] 230[4])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 mux_375_Mux_4_i15_4_lut (.I0(state[2]), .I1(n4943), .I2(state[3]), 
            .I3(state[1]), .O(n1103[4]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_375_Mux_4_i15_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(n63), .I3(n4068), 
            .O(n2106));   // src/timing_controller.v(154[8] 230[4])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i1065_4_lut (.I0(state[3]), .I1(n11356), .I2(n8057), .I3(state[2]), 
            .O(n2144));   // src/timing_controller.v(154[8] 230[4])
    defparam i1065_4_lut.LUT_INIT = 16'h0544;
    SB_DFFSR line_of_data_available_93 (.Q(line_of_data_available), .C(SLM_CLK_c), 
            .D(n2), .R(n6520));   // src/timing_controller.v(88[8] 151[4])
    SB_DFFESR invert_100_i3 (.Q(UPDATE_c_3), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n11506), .R(n4068));   // src/timing_controller.v(160[5] 229[12])
    SB_LUT4 i9964_2_lut (.I0(n4943), .I1(state[3]), .I2(GND_net), .I3(GND_net), 
            .O(n5068));
    defparam i9964_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 sub_71_add_2_27_lut (.I0(GND_net), .I1(state_timeout_counter[25]), 
            .I2(VCC_net), .I3(n10274), .O(n630[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_127 (.I0(fifo_state[2]), .I1(n6461), .I2(fifo_state[0]), 
            .I3(fifo_state[1]), .O(n4_adj_1391));
    defparam i1_2_lut_4_lut_adj_127.LUT_INIT = 16'h00f8;
    SB_LUT4 i12_1_lut_3_lut (.I0(fifo_state[2]), .I1(n6461), .I2(fifo_state[0]), 
            .I3(GND_net), .O(n5));
    defparam i12_1_lut_3_lut.LUT_INIT = 16'h0707;
    SB_LUT4 mux_1004_i1_4_lut (.I0(n11358), .I1(state[1]), .I2(n2144), 
            .I3(n2072), .O(n2145[0]));   // src/timing_controller.v(160[5] 229[12])
    defparam mux_1004_i1_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i1_2_lut_4_lut_adj_128 (.I0(state[1]), .I1(state[2]), .I2(state[0]), 
            .I3(state[3]), .O(n11104));
    defparam i1_2_lut_4_lut_adj_128.LUT_INIT = 16'h0010;
    SB_LUT4 i2_3_lut_4_lut_adj_129 (.I0(state[3]), .I1(n63), .I2(state[1]), 
            .I3(state[2]), .O(n11119));
    defparam i2_3_lut_4_lut_adj_129.LUT_INIT = 16'hffbf;
    
endmodule
//
// Verilog Description of module bluejay_data
//

module bluejay_data (VCC_net, VALID_c, SLM_CLK_c, bluejay_data_out_31__N_920, 
            buffer_switch_done, GND_net, n1459, n3, buffer_switch_done_latched, 
            n5132, n80, n11094, SYNC_c, bluejay_data_out_31__N_919, 
            \state_timeout_counter[7] , line_of_data_available, n5504, 
            n5500, sc32_fifo_almost_empty, n5616, DEBUG_8_c, n106) /* synthesis syn_module_defined=1 */ ;
    input VCC_net;
    output VALID_c;
    input SLM_CLK_c;
    output bluejay_data_out_31__N_920;
    input buffer_switch_done;
    input GND_net;
    output n1459;
    output n3;
    input buffer_switch_done_latched;
    input n5132;
    output n80;
    output n11094;
    output SYNC_c;
    output bluejay_data_out_31__N_919;
    output \state_timeout_counter[7] ;
    input line_of_data_available;
    input n5504;
    input n5500;
    input sc32_fifo_almost_empty;
    input n5616;
    output DEBUG_8_c;
    output n106;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire bluejay_data_out_31__N_921;
    wire [15:0]n963;
    
    wire n5242;
    wire [8:0]n74;
    
    wire n7396, n7403, n5, n4, n147, n5_adj_1384, n11281;
    wire [7:0]state_timeout_counter;   // src/bluejay_data.v(52[11:32])
    
    wire n11285;
    wire [10:0]v_counter_10__N_899;
    wire [10:0]v_counter;   // src/bluejay_data.v(51[12:21])
    
    wire n10322, n109, n5503, n5_adj_1385, n10321, n5_adj_1386;
    wire [3:0]n99;
    
    wire n899, n10380, n6, n11159, n9, n11, n7400, n66, n10320, 
        n10319, n9_adj_1387, n11096, n10686, n10318, n10317, n10316, 
        n10315, n10314, n10313, bluejay_data_out_31__N_918, n10238, 
        n10239, n3464, n1030, n3462, n1026, n3460, n3458, n1017, 
        n11054, n4982, n10244, n10243, n10242, n11279, n12, n7392, 
        n11187, n154, n5470, n5505, n5502, n5501, n11033, n11123, 
        n9351, n10241, n68, n11129, n11038, n10240, n11097, n9_adj_1388, 
        n10538, n10708, n18, n6_adj_1389, n10403;
    
    SB_DFFNESS valid_66 (.Q(VALID_c), .C(SLM_CLK_c), .E(VCC_net), .D(bluejay_data_out_31__N_921), 
            .S(bluejay_data_out_31__N_920));   // src/bluejay_data.v(134[8] 156[4])
    SB_LUT4 i1_2_lut (.I0(n963[9]), .I1(buffer_switch_done), .I2(GND_net), 
            .I3(GND_net), .O(n5242));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 select_621_Select_7_i3_2_lut (.I0(n74[7]), .I1(n1459), .I2(GND_net), 
            .I3(GND_net), .O(n3));   // src/bluejay_data.v(66[9] 129[16])
    defparam select_621_Select_7_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(n963[9]), .I1(n74[7]), .I2(n7396), .I3(n7403), 
            .O(n5));
    defparam i1_4_lut.LUT_INIT = 16'hc0c8;
    SB_LUT4 i1_3_lut (.I0(n1459), .I1(buffer_switch_done_latched), .I2(n74[6]), 
            .I3(GND_net), .O(n4));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i1_2_lut_adj_88 (.I0(n74[6]), .I1(n147), .I2(GND_net), .I3(GND_net), 
            .O(n5_adj_1384));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_88.LUT_INIT = 16'h8888;
    SB_LUT4 i9705_4_lut (.I0(buffer_switch_done_latched), .I1(n963[2]), 
            .I2(n11281), .I3(state_timeout_counter[5]), .O(n11285));
    defparam i9705_4_lut.LUT_INIT = 16'hfefa;
    SB_LUT4 sub_122_add_2_12_lut (.I0(GND_net), .I1(v_counter[10]), .I2(VCC_net), 
            .I3(n10322), .O(v_counter_10__N_899[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4044_4_lut (.I0(n5132), .I1(n1459), .I2(n109), .I3(n74[4]), 
            .O(n5503));   // src/bluejay_data.v(56[8] 131[4])
    defparam i4044_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_2_lut_adj_89 (.I0(n74[4]), .I1(n147), .I2(GND_net), .I3(GND_net), 
            .O(n5_adj_1385));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_89.LUT_INIT = 16'h8888;
    SB_LUT4 sub_122_add_2_11_lut (.I0(GND_net), .I1(v_counter[9]), .I2(VCC_net), 
            .I3(n10321), .O(v_counter_10__N_899[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_90 (.I0(n80), .I1(n147), .I2(GND_net), .I3(GND_net), 
            .O(n5_adj_1386));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_90.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n99[2]), .I1(n74[2]), .I2(n899), .I3(n963[9]), 
            .O(n10380));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2_4_lut.LUT_INIT = 16'hc400;
    SB_CARRY sub_122_add_2_11 (.CI(n10321), .I0(v_counter[9]), .I1(VCC_net), 
            .CO(n10322));
    SB_LUT4 i2_4_lut_adj_91 (.I0(buffer_switch_done_latched), .I1(n10380), 
            .I2(state_timeout_counter[2]), .I3(n963[2]), .O(n6));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2_4_lut_adj_91.LUT_INIT = 16'hfeee;
    SB_LUT4 i3_4_lut (.I0(n74[2]), .I1(n1459), .I2(n963[5]), .I3(n11159), 
            .O(n9));   // src/bluejay_data.v(66[9] 129[16])
    defparam i3_4_lut.LUT_INIT = 16'ha8f8;
    SB_LUT4 i1_2_lut_adj_92 (.I0(n1459), .I1(n7396), .I2(GND_net), .I3(GND_net), 
            .O(n11));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_92.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_93 (.I0(n963[2]), .I1(buffer_switch_done_latched), 
            .I2(GND_net), .I3(GND_net), .O(n11094));
    defparam i1_2_lut_adj_93.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut (.I0(n7400), .I1(n66), .I2(state_timeout_counter[0]), 
            .I3(GND_net), .O(n7403));   // src/bluejay_data.v(56[8] 131[4])
    defparam i2_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 sub_122_add_2_10_lut (.I0(GND_net), .I1(v_counter[8]), .I2(VCC_net), 
            .I3(n10320), .O(v_counter_10__N_899[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_122_add_2_10 (.CI(n10320), .I0(v_counter[8]), .I1(VCC_net), 
            .CO(n10321));
    SB_LUT4 sub_122_add_2_9_lut (.I0(GND_net), .I1(v_counter[7]), .I2(VCC_net), 
            .I3(n10319), .O(v_counter_10__N_899[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_94 (.I0(n963[9]), .I1(n7403), .I2(n74[1]), .I3(GND_net), 
            .O(n9_adj_1387));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_3_lut_adj_94.LUT_INIT = 16'ha8a8;
    SB_CARRY sub_122_add_2_9 (.CI(n10319), .I0(v_counter[7]), .I1(VCC_net), 
            .CO(n10320));
    SB_LUT4 i2_4_lut_adj_95 (.I0(n74[1]), .I1(n11096), .I2(n11), .I3(n9_adj_1387), 
            .O(n10686));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2_4_lut_adj_95.LUT_INIT = 16'hffec;
    SB_DFFESR v_counter_i1 (.Q(v_counter[1]), .C(SLM_CLK_c), .E(n5242), 
            .D(v_counter_10__N_899[1]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i2 (.Q(v_counter[2]), .C(SLM_CLK_c), .E(n5242), 
            .D(v_counter_10__N_899[2]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i3 (.Q(v_counter[3]), .C(SLM_CLK_c), .E(n5242), 
            .D(v_counter_10__N_899[3]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i4 (.Q(v_counter[4]), .C(SLM_CLK_c), .E(n5242), 
            .D(v_counter_10__N_899[4]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i5 (.Q(v_counter[5]), .C(SLM_CLK_c), .E(n5242), 
            .D(v_counter_10__N_899[5]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i6 (.Q(v_counter[6]), .C(SLM_CLK_c), .E(n5242), 
            .D(v_counter_10__N_899[6]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS v_counter_i7 (.Q(v_counter[7]), .C(SLM_CLK_c), .E(n5242), 
            .D(v_counter_10__N_899[7]), .S(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i8 (.Q(v_counter[8]), .C(SLM_CLK_c), .E(n5242), 
            .D(v_counter_10__N_899[8]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i9 (.Q(v_counter[9]), .C(SLM_CLK_c), .E(n5242), 
            .D(v_counter_10__N_899[9]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_LUT4 sub_122_add_2_8_lut (.I0(GND_net), .I1(v_counter[6]), .I2(VCC_net), 
            .I3(n10318), .O(v_counter_10__N_899[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_122_add_2_8 (.CI(n10318), .I0(v_counter[6]), .I1(VCC_net), 
            .CO(n10319));
    SB_LUT4 sub_122_add_2_7_lut (.I0(GND_net), .I1(v_counter[5]), .I2(VCC_net), 
            .I3(n10317), .O(v_counter_10__N_899[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_122_add_2_7 (.CI(n10317), .I0(v_counter[5]), .I1(VCC_net), 
            .CO(n10318));
    SB_DFFESR v_counter_i10 (.Q(v_counter[10]), .C(SLM_CLK_c), .E(n5242), 
            .D(v_counter_10__N_899[10]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_LUT4 sub_122_add_2_6_lut (.I0(GND_net), .I1(v_counter[4]), .I2(VCC_net), 
            .I3(n10316), .O(v_counter_10__N_899[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_122_add_2_6 (.CI(n10316), .I0(v_counter[4]), .I1(VCC_net), 
            .CO(n10317));
    SB_LUT4 sub_122_add_2_5_lut (.I0(GND_net), .I1(v_counter[3]), .I2(VCC_net), 
            .I3(n10315), .O(v_counter_10__N_899[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_122_add_2_5 (.CI(n10315), .I0(v_counter[3]), .I1(VCC_net), 
            .CO(n10316));
    SB_LUT4 sub_122_add_2_4_lut (.I0(GND_net), .I1(v_counter[2]), .I2(VCC_net), 
            .I3(n10314), .O(v_counter_10__N_899[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_122_add_2_4 (.CI(n10314), .I0(v_counter[2]), .I1(VCC_net), 
            .CO(n10315));
    SB_LUT4 sub_122_add_2_3_lut (.I0(GND_net), .I1(v_counter[1]), .I2(VCC_net), 
            .I3(n10313), .O(v_counter_10__N_899[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_122_add_2_3 (.CI(n10313), .I0(v_counter[1]), .I1(VCC_net), 
            .CO(n10314));
    SB_LUT4 sub_122_add_2_2_lut (.I0(GND_net), .I1(v_counter[0]), .I2(n899), 
            .I3(VCC_net), .O(v_counter_10__N_899[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_122_add_2_2 (.CI(VCC_net), .I0(v_counter[0]), .I1(n899), 
            .CO(n10313));
    SB_DFFN sync_68 (.Q(SYNC_c), .C(SLM_CLK_c), .D(bluejay_data_out_31__N_918));   // src/bluejay_data.v(134[8] 156[4])
    SB_LUT4 sub_120_add_2_3_lut (.I0(GND_net), .I1(state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n10238), .O(n74[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_120_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_120_add_2_3 (.CI(n10238), .I0(state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n10239));
    SB_DFFSR state_FSM_i10 (.Q(n963[9]), .C(SLM_CLK_c), .D(n3464), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i9 (.Q(bluejay_data_out_31__N_921), .C(SLM_CLK_c), 
            .D(n1030), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_LUT4 sub_120_add_2_2_lut (.I0(GND_net), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n74[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_120_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR state_FSM_i8 (.Q(bluejay_data_out_31__N_920), .C(SLM_CLK_c), 
            .D(n3462), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i7 (.Q(bluejay_data_out_31__N_919), .C(SLM_CLK_c), 
            .D(n1026), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i6 (.Q(n963[5]), .C(SLM_CLK_c), .D(n3460), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i5 (.Q(n963[4]), .C(SLM_CLK_c), .D(n3458), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i4 (.Q(bluejay_data_out_31__N_918), .C(SLM_CLK_c), 
            .D(n1017), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i3 (.Q(n963[2]), .C(SLM_CLK_c), .D(n11054), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i2 (.Q(n963[1]), .C(SLM_CLK_c), .D(n4982), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_CARRY sub_120_add_2_2 (.CI(VCC_net), .I0(state_timeout_counter[0]), 
            .I1(GND_net), .CO(n10238));
    SB_LUT4 sub_120_add_2_9_lut (.I0(GND_net), .I1(\state_timeout_counter[7] ), 
            .I2(VCC_net), .I3(n10244), .O(n74[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_120_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_120_add_2_8_lut (.I0(GND_net), .I1(state_timeout_counter[6]), 
            .I2(VCC_net), .I3(n10243), .O(n74[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_120_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_120_add_2_8 (.CI(n10243), .I0(state_timeout_counter[6]), 
            .I1(VCC_net), .CO(n10244));
    SB_LUT4 sub_120_add_2_7_lut (.I0(n11279), .I1(state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n10242), .O(n11281)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_120_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_120_add_2_7 (.CI(n10242), .I0(state_timeout_counter[5]), 
            .I1(VCC_net), .CO(n10243));
    SB_LUT4 i1_2_lut_adj_96 (.I0(line_of_data_available), .I1(n12), .I2(GND_net), 
            .I3(GND_net), .O(n7392));   // src/top.v(468[6:28])
    defparam i1_2_lut_adj_96.LUT_INIT = 16'heeee;
    SB_LUT4 i9611_4_lut (.I0(n963[5]), .I1(n66), .I2(state_timeout_counter[0]), 
            .I3(n7392), .O(n11187));
    defparam i9611_4_lut.LUT_INIT = 16'haa8a;
    SB_LUT4 i140_4_lut (.I0(n11187), .I1(n7400), .I2(n963[9]), .I3(n154), 
            .O(n147));   // src/bluejay_data.v(66[9] 129[16])
    defparam i140_4_lut.LUT_INIT = 16'hfaba;
    SB_LUT4 i2_3_lut_adj_97 (.I0(bluejay_data_out_31__N_920), .I1(n963[4]), 
            .I2(n963[1]), .I3(GND_net), .O(n1459));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2_3_lut_adj_97.LUT_INIT = 16'hfefe;
    SB_LUT4 i9699_2_lut (.I0(n1459), .I1(n147), .I2(GND_net), .I3(GND_net), 
            .O(n11279));
    defparam i9699_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESS state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(SLM_CLK_c), 
            .E(n5132), .D(n10686), .S(n5470));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(SLM_CLK_c), 
            .E(n5132), .D(n9), .S(n5505));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(SLM_CLK_c), 
            .E(n5132), .D(n5_adj_1386), .S(n5504));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(SLM_CLK_c), 
            .E(n5132), .D(n5_adj_1385), .S(n5503));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS state_timeout_counter_i0_i5 (.Q(state_timeout_counter[5]), .C(SLM_CLK_c), 
            .E(n5132), .D(n11285), .S(n5502));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS state_timeout_counter_i0_i6 (.Q(state_timeout_counter[6]), .C(SLM_CLK_c), 
            .E(n5132), .D(n5_adj_1384), .S(n5501));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS state_timeout_counter_i0_i7 (.Q(\state_timeout_counter[7] ), 
            .C(SLM_CLK_c), .E(n5132), .D(n5), .S(n5500));   // src/bluejay_data.v(56[8] 131[4])
    SB_LUT4 i2_3_lut_4_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[5]), 
            .I2(n66), .I3(n11033), .O(n11123));   // src/bluejay_data.v(56[8] 131[4])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[5]), 
            .I2(n9351), .I3(GND_net), .O(n12));   // src/bluejay_data.v(56[8] 131[4])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_98 (.I0(state_timeout_counter[0]), .I1(state_timeout_counter[4]), 
            .I2(state_timeout_counter[3]), .I3(GND_net), .O(n154));
    defparam i1_2_lut_3_lut_adj_98.LUT_INIT = 16'hfdfd;
    SB_LUT4 sub_120_add_2_6_lut (.I0(GND_net), .I1(state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n10241), .O(n74[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_120_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i349_2_lut_3_lut_4_lut (.I0(n154), .I1(n12), .I2(line_of_data_available), 
            .I3(n963[1]), .O(n1017));   // src/bluejay_data.v(69[17] 76[20])
    defparam i349_2_lut_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_CARRY sub_120_add_2_6 (.CI(n10241), .I0(state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n10242));
    SB_LUT4 i362_2_lut_4_lut (.I0(n154), .I1(n12), .I2(sc32_fifo_almost_empty), 
            .I3(bluejay_data_out_31__N_920), .O(n1030));   // src/bluejay_data.v(66[9] 129[16])
    defparam i362_2_lut_4_lut.LUT_INIT = 16'hf100;
    SB_LUT4 i19_2_lut_3_lut (.I0(n154), .I1(n12), .I2(sc32_fifo_almost_empty), 
            .I3(GND_net), .O(n68));   // src/bluejay_data.v(97[21:87])
    defparam i19_2_lut_3_lut.LUT_INIT = 16'hf1f1;
    SB_LUT4 i1_2_lut_4_lut (.I0(n11129), .I1(\state_timeout_counter[7] ), 
            .I2(state_timeout_counter[6]), .I3(state_timeout_counter[2]), 
            .O(n11038));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9583_2_lut_3_lut (.I0(line_of_data_available), .I1(n154), .I2(n12), 
            .I3(GND_net), .O(n11159));
    defparam i9583_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 sub_120_add_2_5_lut (.I0(GND_net), .I1(state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n10240), .O(n80)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_120_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_99 (.I0(state_timeout_counter[0]), .I1(n963[2]), 
            .I2(buffer_switch_done_latched), .I3(GND_net), .O(n11097));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_3_lut_adj_99.LUT_INIT = 16'h0808;
    SB_DFFN get_next_word_67 (.Q(DEBUG_8_c), .C(SLM_CLK_c), .D(n5616));   // src/bluejay_data.v(134[8] 156[4])
    SB_LUT4 i1_3_lut_4_lut (.I0(buffer_switch_done_latched), .I1(n963[1]), 
            .I2(n154), .I3(n12), .O(n4982));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'heeea;
    SB_LUT4 i1_3_lut_adj_100 (.I0(n963[9]), .I1(n7403), .I2(n74[0]), .I3(GND_net), 
            .O(n9_adj_1388));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_3_lut_adj_100.LUT_INIT = 16'ha8a8;
    SB_LUT4 i2_4_lut_adj_101 (.I0(n11123), .I1(n963[9]), .I2(n11038), 
            .I3(state_timeout_counter[0]), .O(n10538));
    defparam i2_4_lut_adj_101.LUT_INIT = 16'h0400;
    SB_LUT4 i1_4_lut_adj_102 (.I0(n963[2]), .I1(n10538), .I2(n963[1]), 
            .I3(n11159), .O(n11054));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_4_lut_adj_102.LUT_INIT = 16'heefe;
    SB_CARRY sub_120_add_2_5 (.CI(n10240), .I0(state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n10241));
    SB_LUT4 i2_4_lut_adj_103 (.I0(n74[0]), .I1(n11097), .I2(n11), .I3(n9_adj_1388), 
            .O(n10708));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2_4_lut_adj_103.LUT_INIT = 16'hffec;
    SB_LUT4 equal_123_i18_2_lut (.I0(v_counter[9]), .I1(v_counter[10]), 
            .I2(GND_net), .I3(GND_net), .O(n18));   // src/bluejay_data.v(109[25:41])
    defparam equal_123_i18_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_104 (.I0(v_counter[2]), .I1(v_counter[3]), .I2(v_counter[4]), 
            .I3(v_counter[5]), .O(n6_adj_1389));
    defparam i2_4_lut_adj_104.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_105 (.I0(v_counter[0]), .I1(n6_adj_1389), .I2(n18), 
            .I3(v_counter[1]), .O(n11129));
    defparam i3_4_lut_adj_105.LUT_INIT = 16'hfffd;
    SB_LUT4 i2_3_lut_adj_106 (.I0(v_counter[7]), .I1(v_counter[8]), .I2(v_counter[6]), 
            .I3(GND_net), .O(n11033));   // src/bluejay_data.v(56[8] 131[4])
    defparam i2_3_lut_adj_106.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_107 (.I0(n11033), .I1(n11129), .I2(GND_net), 
            .I3(GND_net), .O(n99[2]));   // src/bluejay_data.v(56[8] 131[4])
    defparam i1_2_lut_adj_107.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_108 (.I0(buffer_switch_done_latched), .I1(line_of_data_available), 
            .I2(n963[5]), .I3(n899), .O(n10403));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2_4_lut_adj_108.LUT_INIT = 16'h5010;
    SB_LUT4 i2014_4_lut (.I0(n10403), .I1(n963[9]), .I2(n99[2]), .I3(n899), 
            .O(n3460));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2014_4_lut.LUT_INIT = 16'haaea;
    SB_LUT4 sub_120_add_2_4_lut (.I0(GND_net), .I1(state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n10239), .O(n74[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_120_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2016_4_lut (.I0(buffer_switch_done_latched), .I1(bluejay_data_out_31__N_919), 
            .I2(n68), .I3(bluejay_data_out_31__N_920), .O(n3462));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2016_4_lut.LUT_INIT = 16'hcdcc;
    SB_LUT4 i2018_3_lut_4_lut (.I0(buffer_switch_done_latched), .I1(n899), 
            .I2(bluejay_data_out_31__N_921), .I3(n963[9]), .O(n3464));   // src/bluejay_data.v(62[9] 65[12])
    defparam i2018_3_lut_4_lut.LUT_INIT = 16'hf4f0;
    SB_LUT4 i2012_3_lut_4_lut (.I0(buffer_switch_done_latched), .I1(n899), 
            .I2(bluejay_data_out_31__N_918), .I3(n963[4]), .O(n3458));   // src/bluejay_data.v(62[9] 65[12])
    defparam i2012_3_lut_4_lut.LUT_INIT = 16'hf4f0;
    SB_DFFESS state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(SLM_CLK_c), 
            .E(n5132), .D(n10708), .S(n5470));   // src/bluejay_data.v(56[8] 131[4])
    SB_LUT4 i1_2_lut_3_lut_adj_109 (.I0(n11033), .I1(n11129), .I2(n12), 
            .I3(GND_net), .O(n7400));   // src/bluejay_data.v(109[25:41])
    defparam i1_2_lut_3_lut_adj_109.LUT_INIT = 16'h0e0e;
    SB_CARRY sub_120_add_2_4 (.CI(n10239), .I0(state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n10240));
    SB_DFFESR v_counter_i0 (.Q(v_counter[0]), .C(SLM_CLK_c), .E(n5242), 
            .D(v_counter_10__N_899[0]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_LUT4 reduce_or_357_i1_4_lut_4_lut (.I0(n899), .I1(line_of_data_available), 
            .I2(n963[4]), .I3(n963[5]), .O(n1026));   // src/bluejay_data.v(69[17] 76[20])
    defparam reduce_or_357_i1_4_lut_4_lut.LUT_INIT = 16'h5450;
    SB_LUT4 i1_2_lut_3_lut_adj_110 (.I0(state_timeout_counter[1]), .I1(n963[2]), 
            .I2(buffer_switch_done_latched), .I3(GND_net), .O(n11096));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_3_lut_adj_110.LUT_INIT = 16'h0808;
    SB_LUT4 i4011_3_lut_3_lut (.I0(buffer_switch_done), .I1(bluejay_data_out_31__N_919), 
            .I2(bluejay_data_out_31__N_918), .I3(GND_net), .O(n5470));   // src/bluejay_data.v(56[8] 131[4])
    defparam i4011_3_lut_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_3_lut_4_lut_adj_111 (.I0(n963[5]), .I1(state_timeout_counter[0]), 
            .I2(n66), .I3(n7392), .O(n7396));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_3_lut_4_lut_adj_111.LUT_INIT = 16'haaa2;
    SB_LUT4 i4046_4_lut_4_lut (.I0(buffer_switch_done), .I1(bluejay_data_out_31__N_921), 
            .I2(n6), .I3(bluejay_data_out_31__N_919), .O(n5505));   // src/bluejay_data.v(56[8] 131[4])
    defparam i4046_4_lut_4_lut.LUT_INIT = 16'h5554;
    SB_LUT4 i1_2_lut_3_lut_adj_112 (.I0(state_timeout_counter[3]), .I1(n963[2]), 
            .I2(buffer_switch_done_latched), .I3(GND_net), .O(n106));   // src/bluejay_data.v(62[9] 65[12])
    defparam i1_2_lut_3_lut_adj_112.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_3_lut_adj_113 (.I0(state_timeout_counter[4]), .I1(n963[2]), 
            .I2(buffer_switch_done_latched), .I3(GND_net), .O(n109));   // src/bluejay_data.v(62[9] 65[12])
    defparam i1_2_lut_3_lut_adj_113.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_adj_114 (.I0(state_timeout_counter[4]), .I1(state_timeout_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n66));
    defparam i1_2_lut_adj_114.LUT_INIT = 16'heeee;
    SB_LUT4 i4043_2_lut_2_lut (.I0(buffer_switch_done), .I1(bluejay_data_out_31__N_919), 
            .I2(GND_net), .I3(GND_net), .O(n5502));   // src/bluejay_data.v(56[8] 131[4])
    defparam i4043_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_3_lut_adj_115 (.I0(\state_timeout_counter[7] ), .I1(state_timeout_counter[6]), 
            .I2(state_timeout_counter[2]), .I3(GND_net), .O(n9351));   // src/bluejay_data.v(56[8] 131[4])
    defparam i2_3_lut_adj_115.LUT_INIT = 16'hfefe;
    SB_LUT4 i4042_4_lut_4_lut (.I0(buffer_switch_done), .I1(n963[2]), .I2(n4), 
            .I3(state_timeout_counter[6]), .O(n5501));   // src/bluejay_data.v(56[8] 131[4])
    defparam i4042_4_lut_4_lut.LUT_INIT = 16'h5450;
    SB_LUT4 i1_2_lut_adj_116 (.I0(n154), .I1(n12), .I2(GND_net), .I3(GND_net), 
            .O(n899));   // src/bluejay_data.v(56[8] 131[4])
    defparam i1_2_lut_adj_116.LUT_INIT = 16'heeee;
    
endmodule
//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=20) 
//

module \uart_rx(CLKS_PER_BIT=20)  (SLM_CLK_c, r_SM_Main, \r_SM_Main_2__N_949[2] , 
            GND_net, n8012, r_Rx_Data, n5214, n4, n5709, pc_data_rx, 
            n5692, n5527, n4_adj_1, UART_RX_c, n5665, n5658, n5656, 
            n4_adj_2, \r_Bit_Index[0] , n6690, n5644, n5643, n5825, 
            n10608, VCC_net, debug_led3, n5821, n5019) /* synthesis syn_module_defined=1 */ ;
    input SLM_CLK_c;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_949[2] ;
    input GND_net;
    output n8012;
    output r_Rx_Data;
    output n5214;
    output n4;
    input n5709;
    output [7:0]pc_data_rx;
    input n5692;
    output n5527;
    output n4_adj_1;
    input UART_RX_c;
    input n5665;
    input n5658;
    input n5656;
    output n4_adj_2;
    output \r_Bit_Index[0] ;
    output n6690;
    input n5644;
    input n5643;
    input n5825;
    input n10608;
    input VCC_net;
    output debug_led3;
    input n5821;
    output n5019;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [9:0]n45;
    
    wire n6719;
    wire [9:0]r_Clock_Count;   // src/uart_rx.v(32[17:30])
    
    wire n6711, n11173;
    wire [2:0]r_Bit_Index;   // src/uart_rx.v(33[17:28])
    
    wire n116, n6, n3, r_Rx_Data_R;
    wire [2:0]n340;
    
    wire n126, n6752, n119, n10340, n10339, n10338, n6705, n10690, 
        n10337, n122, n10336, n10335, n10334, n10333, n10332, 
        n10442, n111, n6_adj_1383, n8, n11253;
    
    SB_DFFESR r_Clock_Count_1349__i0 (.Q(r_Clock_Count[0]), .C(SLM_CLK_c), 
            .E(n6719), .D(n45[0]), .R(n6711));   // src/uart_rx.v(120[34:51])
    SB_LUT4 i9597_2_lut (.I0(r_SM_Main[1]), .I1(\r_SM_Main_2__N_949[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n11173));
    defparam i9597_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6566_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8012));
    defparam i6566_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut (.I0(n116), .I1(r_SM_Main[1]), .I2(GND_net), .I3(GND_net), 
            .O(n6));   // src/uart_rx.v(36[17:26])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(SLM_CLK_c), .D(n3), .R(r_SM_Main[2]));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(SLM_CLK_c), .D(r_Rx_Data_R));   // src/uart_rx.v(41[10] 45[8])
    SB_LUT4 i1_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[2]), .I2(n6), .I3(r_SM_Main[0]), 
            .O(n6719));   // src/uart_rx.v(36[17:26])
    defparam i1_4_lut.LUT_INIT = 16'h3133;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(\r_SM_Main_2__N_949[2] ), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main[2]), .O(n5214));   // src/uart_rx.v(49[10] 144[8])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h000d;
    SB_LUT4 equal_149_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // src/uart_rx.v(97[17:39])
    defparam equal_149_i4_2_lut.LUT_INIT = 16'heeee;
    SB_DFF r_Rx_Byte_i7 (.Q(pc_data_rx[7]), .C(SLM_CLK_c), .D(n5709));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(pc_data_rx[6]), .C(SLM_CLK_c), .D(n5692));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(SLM_CLK_c), .E(n5214), 
            .D(n340[1]), .R(n5527));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 equal_147_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // src/uart_rx.v(97[17:39])
    defparam equal_147_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(SLM_CLK_c), .D(UART_RX_c));   // src/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Byte_i5 (.Q(pc_data_rx[5]), .C(SLM_CLK_c), .D(n5665));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(SLM_CLK_c), .E(n5214), 
            .D(n340[2]), .R(n5527));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i5296_3_lut (.I0(r_SM_Main[1]), .I1(n126), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n6752));   // src/uart_rx.v(36[17:26])
    defparam i5296_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(SLM_CLK_c), .D(n6752), 
            .R(r_SM_Main[2]));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(pc_data_rx[4]), .C(SLM_CLK_c), .D(n5658));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(pc_data_rx[3]), .C(SLM_CLK_c), .D(n5656));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 equal_144_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // src/uart_rx.v(97[17:39])
    defparam equal_144_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i4068_3_lut (.I0(n5214), .I1(r_SM_Main[1]), .I2(n119), .I3(GND_net), 
            .O(n5527));   // src/uart_rx.v(49[10] 144[8])
    defparam i4068_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 i2_3_lut_4_lut_adj_85 (.I0(r_SM_Main[2]), .I1(n11173), .I2(r_SM_Main[0]), 
            .I3(\r_Bit_Index[0] ), .O(n6690));   // src/uart_rx.v(49[10] 144[8])
    defparam i2_3_lut_4_lut_adj_85.LUT_INIT = 16'h0400;
    SB_LUT4 i1510_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n340[1]));   // src/uart_rx.v(102[36:51])
    defparam i1510_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 r_Clock_Count_1349_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[9]), .I3(n10340), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1349_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1349_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n10339), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1349_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1349_add_4_10 (.CI(n10339), .I0(GND_net), .I1(r_Clock_Count[8]), 
            .CO(n10340));
    SB_DFF r_Rx_Byte_i2 (.Q(pc_data_rx[2]), .C(SLM_CLK_c), .D(n5644));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(pc_data_rx[1]), .C(SLM_CLK_c), .D(n5643));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_Clock_Count_1349_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n10338), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1349_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1349_add_4_9 (.CI(n10338), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n10339));
    SB_DFF r_Rx_Byte_i0 (.Q(pc_data_rx[0]), .C(SLM_CLK_c), .D(n5825));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Rx_DV_52 (.Q(debug_led3), .C(SLM_CLK_c), .E(VCC_net), .D(n10608));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i5249_3_lut (.I0(n116), .I1(\r_SM_Main_2__N_949[2] ), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n6705));   // src/uart_rx.v(36[17:26])
    defparam i5249_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i12_4_lut (.I0(r_Rx_Data), .I1(n119), .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_949[2] ), 
            .O(n10690));   // src/uart_rx.v(30[17:26])
    defparam i12_4_lut.LUT_INIT = 16'hc505;
    SB_LUT4 i5284_3_lut (.I0(n10690), .I1(n6705), .I2(r_SM_Main[0]), .I3(GND_net), 
            .O(n3));   // src/uart_rx.v(36[17:26])
    defparam i5284_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 r_Clock_Count_1349_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n10337), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1349_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1349_add_4_8 (.CI(n10337), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n10338));
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(SLM_CLK_c), .D(n122));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_Clock_Count_1349_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n10336), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1349_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1349_add_4_7 (.CI(n10336), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n10337));
    SB_LUT4 r_Clock_Count_1349_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n10335), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1349_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1349_add_4_6 (.CI(n10335), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n10336));
    SB_LUT4 r_Clock_Count_1349_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n10334), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1349_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1349_add_4_5 (.CI(n10334), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n10335));
    SB_LUT4 r_Clock_Count_1349_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n10333), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1349_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1349_add_4_4 (.CI(n10333), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n10334));
    SB_LUT4 r_Clock_Count_1349_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n10332), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1349_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1349_add_4_3 (.CI(n10332), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n10333));
    SB_DFFESR r_Clock_Count_1349__i1 (.Q(r_Clock_Count[1]), .C(SLM_CLK_c), 
            .E(n6719), .D(n45[1]), .R(n6711));   // src/uart_rx.v(120[34:51])
    SB_DFFE r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n5821));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_Clock_Count_1349_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1349_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Clock_Count_1349__i2 (.Q(r_Clock_Count[2]), .C(SLM_CLK_c), 
            .E(n6719), .D(n45[2]), .R(n6711));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1349__i3 (.Q(r_Clock_Count[3]), .C(SLM_CLK_c), 
            .E(n6719), .D(n45[3]), .R(n6711));   // src/uart_rx.v(120[34:51])
    SB_CARRY r_Clock_Count_1349_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n10332));
    SB_DFFESR r_Clock_Count_1349__i4 (.Q(r_Clock_Count[4]), .C(SLM_CLK_c), 
            .E(n6719), .D(n45[4]), .R(n6711));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1349__i5 (.Q(r_Clock_Count[5]), .C(SLM_CLK_c), 
            .E(n6719), .D(n45[5]), .R(n6711));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1349__i6 (.Q(r_Clock_Count[6]), .C(SLM_CLK_c), 
            .E(n6719), .D(n45[6]), .R(n6711));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1349__i7 (.Q(r_Clock_Count[7]), .C(SLM_CLK_c), 
            .E(n6719), .D(n45[7]), .R(n6711));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1349__i8 (.Q(r_Clock_Count[8]), .C(SLM_CLK_c), 
            .E(n6719), .D(n45[8]), .R(n6711));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1349__i9 (.Q(r_Clock_Count[9]), .C(SLM_CLK_c), 
            .E(n6719), .D(n45[9]), .R(n6711));   // src/uart_rx.v(120[34:51])
    SB_LUT4 i2_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[2]), .O(n10442));   // src/uart_rx.v(32[17:30])
    defparam i2_4_lut.LUT_INIT = 16'hffec;
    SB_LUT4 i1_3_lut (.I0(n111), .I1(r_Clock_Count[4]), .I2(n10442), .I3(GND_net), 
            .O(\r_SM_Main_2__N_949[2] ));   // src/uart_rx.v(32[17:30])
    defparam i1_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[9]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_1383));   // src/uart_rx.v(32[17:30])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[7]), .I2(r_Clock_Count[5]), 
            .I3(n6_adj_1383), .O(n111));   // src/uart_rx.v(32[17:30])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[4]), .I2(r_Clock_Count[0]), 
            .I3(n111), .O(n8));
    defparam i3_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i4_3_lut (.I0(r_Clock_Count[1]), .I1(n8), .I2(r_Clock_Count[2]), 
            .I3(GND_net), .O(n116));
    defparam i4_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9675_3_lut (.I0(r_SM_Main[0]), .I1(n116), .I2(r_Rx_Data), 
            .I3(GND_net), .O(n11253));
    defparam i9675_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i5295_3_lut_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(\r_SM_Main_2__N_949[2] ), 
            .I2(r_Rx_Data), .I3(n116), .O(n126));   // src/uart_rx.v(49[10] 144[8])
    defparam i5295_3_lut_4_lut_4_lut.LUT_INIT = 16'hddd8;
    SB_LUT4 i1_4_lut_adj_86 (.I0(r_SM_Main[2]), .I1(n11253), .I2(\r_SM_Main_2__N_949[2] ), 
            .I3(r_SM_Main[1]), .O(n6711));   // src/uart_rx.v(36[17:26])
    defparam i1_4_lut_adj_86.LUT_INIT = 16'h5011;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), 
            .I2(\r_SM_Main_2__N_949[2] ), .I3(r_SM_Main[0]), .O(n122));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i1517_2_lut_3_lut (.I0(\r_Bit_Index[0] ), .I1(r_Bit_Index[1]), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n340[2]));   // src/uart_rx.v(49[10] 144[8])
    defparam i1517_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i4_4_lut_adj_87 (.I0(\r_Bit_Index[0] ), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(n11173), .O(n5019));   // src/uart_rx.v(49[10] 144[8])
    defparam i4_4_lut_adj_87.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_2_lut_3_lut (.I0(\r_Bit_Index[0] ), .I1(r_Bit_Index[1]), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n119));   // src/uart_rx.v(49[10] 144[8])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    
endmodule
//
// Verilog Description of module clock
//

module clock (GND_net, VCC_net, ICE_SYSCLK_c, pll_clk_unbuf) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    input ICE_SYSCLK_c;
    output pll_clk_unbuf;
    
    
    SB_PLL40_CORE pll_config (.REFERENCECLK(ICE_SYSCLK_c), .PLLOUTGLOBAL(pll_clk_unbuf), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=15, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=222, LSE_RLINE=228 */ ;   // src/top.v(222[7] 228[3])
    defparam pll_config.FEEDBACK_PATH = "SIMPLE";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll_config.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll_config.FDA_FEEDBACK = 0;
    defparam pll_config.FDA_RELATIVE = 0;
    defparam pll_config.PLLOUT_SELECT = "GENCLK";
    defparam pll_config.DIVR = 4'b0001;
    defparam pll_config.DIVF = 7'b1010010;
    defparam pll_config.DIVQ = 3'b100;
    defparam pll_config.FILTER_RANGE = 3'b001;
    defparam pll_config.ENABLE_ICEGATE = 1'b0;
    defparam pll_config.TEST_MODE = 1'b0;
    defparam pll_config.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module spi
//

module spi (VCC_net, GND_net, SLM_CLK_c, SEN_c_1, SOUT_c, n5113, 
            \rx_shift_reg[0] , n2329, multi_byte_spi_trans_flag_r, spi_start_transfer_r, 
            tx_addr_byte, n5081, SDAT_c_15, n5706, \rx_shift_reg[1] , 
            n5705, \rx_shift_reg[2] , n5704, \rx_shift_reg[3] , n5703, 
            \rx_shift_reg[4] , n5702, \rx_shift_reg[5] , n5701, \rx_shift_reg[6] , 
            n5700, \rx_shift_reg[7] , n5699, rx_buf_byte, n5698, n5697, 
            n5696, n5695, n5694, \tx_data_byte[1] , \tx_shift_reg[0] , 
            \tx_data_byte[2] , \tx_data_byte[3] , \tx_data_byte[4] , n5693, 
            \tx_data_byte[5] , \tx_data_byte[6] , \tx_data_byte[7] , spi_rx_byte_ready, 
            SCK_c_0, n5120, n10792, n5621) /* synthesis syn_module_defined=1 */ ;
    input VCC_net;
    input GND_net;
    input SLM_CLK_c;
    output SEN_c_1;
    input SOUT_c;
    output n5113;
    output \rx_shift_reg[0] ;
    output n2329;
    input multi_byte_spi_trans_flag_r;
    input spi_start_transfer_r;
    input [7:0]tx_addr_byte;
    output n5081;
    output SDAT_c_15;
    input n5706;
    output \rx_shift_reg[1] ;
    input n5705;
    output \rx_shift_reg[2] ;
    input n5704;
    output \rx_shift_reg[3] ;
    input n5703;
    output \rx_shift_reg[4] ;
    input n5702;
    output \rx_shift_reg[5] ;
    input n5701;
    output \rx_shift_reg[6] ;
    input n5700;
    output \rx_shift_reg[7] ;
    input n5699;
    output [7:0]rx_buf_byte;
    input n5698;
    input n5697;
    input n5696;
    input n5695;
    input n5694;
    input \tx_data_byte[1] ;
    output \tx_shift_reg[0] ;
    input \tx_data_byte[2] ;
    input \tx_data_byte[3] ;
    input \tx_data_byte[4] ;
    input n5693;
    input \tx_data_byte[5] ;
    input \tx_data_byte[6] ;
    input \tx_data_byte[7] ;
    output spi_rx_byte_ready;
    output SCK_c_0;
    output n5120;
    input n10792;
    input n5621;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [9:0]n45;
    wire [9:0]counter;   // src/spi.v(69[11:18])
    
    wire n10328;
    wire [7:0]n2406;
    wire [3:0]state;   // src/spi.v(71[11:16])
    
    wire n11372, n10329, n5142, n5487, n19, n11407, n11247, n37, 
        n14, n35, n10327;
    wire [2:0]n1105;
    
    wire n10326, n10325;
    wire [3:0]state_3__N_1122;
    
    wire n11090, n10324, n10323, n5012, n4, n11277, n11039, n11418, 
        n3, n16, n24;
    wire [15:0]tx_shift_reg;   // src/spi.v(70[12:24])
    wire [15:0]n2330;
    
    wire n3_adj_1373, n21;
    wire [7:0]n315;
    wire [7:0]multi_byte_counter;   // src/spi.v(68[11:29])
    
    wire n10312, n10311, n10310, n5199, n5517, n11370, n5009, 
        n10309, n19_adj_1374, n11091, n5179, n10308, n5171, n5172, 
        n11416, n11030, n7, n11089, n3_adj_1375, n11237, n4_adj_1376, 
        n22, n11273, n4813, n10307, n11366, n7_adj_1377, n10306, 
        n8, n10331, n10330, n11397, n11398, n14_adj_1378, n10, 
        n4931, n10_adj_1379, n14_adj_1380;
    
    SB_LUT4 counter_1347_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[6]), 
            .I3(n10328), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1347_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9850_2_lut (.I0(n2406[6]), .I1(state[3]), .I2(GND_net), .I3(GND_net), 
            .O(n11372));
    defparam i9850_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1347_add_4_8 (.CI(n10328), .I0(VCC_net), .I1(counter[6]), 
            .CO(n10329));
    SB_DFFESR counter_1347__i0 (.Q(counter[0]), .C(SLM_CLK_c), .E(n5142), 
            .D(n45[0]), .R(n5487));   // src/spi.v(183[28:41])
    SB_LUT4 i9858_3_lut (.I0(state[0]), .I1(state[2]), .I2(n19), .I3(GND_net), 
            .O(n11407));
    defparam i9858_3_lut.LUT_INIT = 16'h4d4d;
    SB_LUT4 i66_4_lut (.I0(n11247), .I1(n11372), .I2(state[1]), .I3(state[2]), 
            .O(n37));
    defparam i66_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i1_4_lut (.I0(state[3]), .I1(n14), .I2(n11407), .I3(state[1]), 
            .O(n35));
    defparam i1_4_lut.LUT_INIT = 16'h5011;
    SB_LUT4 i1_4_lut_adj_69 (.I0(n35), .I1(n37), .I2(state[0]), .I3(state[2]), 
            .O(n5487));
    defparam i1_4_lut_adj_69.LUT_INIT = 16'haaae;
    SB_LUT4 counter_1347_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[5]), 
            .I3(n10327), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1347_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF byte_recv_92_i2 (.Q(SEN_c_1), .C(SLM_CLK_c), .D(n1105[1]));   // src/spi.v(88[9] 219[16])
    SB_CARRY counter_1347_add_4_7 (.CI(n10327), .I0(VCC_net), .I1(counter[5]), 
            .CO(n10328));
    SB_LUT4 counter_1347_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[4]), 
            .I3(n10326), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1347_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1347_add_4_6 (.CI(n10326), .I0(VCC_net), .I1(counter[4]), 
            .CO(n10327));
    SB_DFFE rx_shift_reg_i0 (.Q(\rx_shift_reg[0] ), .C(SLM_CLK_c), .E(n5113), 
            .D(SOUT_c));   // src/spi.v(76[8] 221[4])
    SB_LUT4 counter_1347_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[3]), 
            .I3(n10325), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1347_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFE state_i0 (.Q(state[0]), .C(SLM_CLK_c), .E(n11090), .D(state_3__N_1122[0]));   // src/spi.v(76[8] 221[4])
    SB_CARRY counter_1347_add_4_5 (.CI(n10325), .I0(VCC_net), .I1(counter[3]), 
            .CO(n10326));
    SB_LUT4 counter_1347_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[2]), 
            .I3(n10324), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1347_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1347_add_4_4 (.CI(n10324), .I0(VCC_net), .I1(counter[2]), 
            .CO(n10325));
    SB_LUT4 counter_1347_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[1]), 
            .I3(n10323), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1347_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9992_4_lut (.I0(state[3]), .I1(state[1]), .I2(n5012), .I3(n14), 
            .O(n5142));   // src/spi.v(88[9] 219[16])
    defparam i9992_4_lut.LUT_INIT = 16'h4c5f;
    SB_LUT4 i1_4_lut_adj_70 (.I0(state[0]), .I1(state[1]), .I2(state[3]), 
            .I3(state[2]), .O(n4));
    defparam i1_4_lut_adj_70.LUT_INIT = 16'h081c;
    SB_LUT4 i9685_2_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(state[2]), 
            .I3(GND_net), .O(n11277));   // src/spi.v(88[9] 219[16])
    defparam i9685_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i1_3_lut (.I0(counter[4]), .I1(n4), .I2(n11039), .I3(GND_net), 
            .O(n2329));
    defparam i1_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i9890_2_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(state[2]), 
            .I3(GND_net), .O(n11418));   // src/spi.v(88[9] 219[16])
    defparam i9890_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_CARRY counter_1347_add_4_3 (.CI(n10323), .I0(VCC_net), .I1(counter[1]), 
            .CO(n10324));
    SB_LUT4 mux_56_Mux_1_i3_3_lut_3_lut (.I0(multi_byte_spi_trans_flag_r), 
            .I1(state[0]), .I2(state[1]), .I3(GND_net), .O(n3));
    defparam mux_56_Mux_1_i3_3_lut_3_lut.LUT_INIT = 16'h3e3e;
    SB_LUT4 i1_4_lut_adj_71 (.I0(n11039), .I1(state[3]), .I2(counter[4]), 
            .I3(state[1]), .O(n16));   // src/spi.v(88[9] 219[16])
    defparam i1_4_lut_adj_71.LUT_INIT = 16'hf5c4;
    SB_LUT4 i30_4_lut (.I0(spi_start_transfer_r), .I1(state[3]), .I2(state[1]), 
            .I3(state[0]), .O(n24));   // src/spi.v(88[9] 219[16])
    defparam i30_4_lut.LUT_INIT = 16'hcfc1;
    SB_LUT4 mux_1117_i16_3_lut (.I0(tx_addr_byte[7]), .I1(tx_shift_reg[14]), 
            .I2(n2329), .I3(GND_net), .O(n2330[15]));   // src/spi.v(88[9] 219[16])
    defparam mux_1117_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_1347_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1347_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1347_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n10323));
    SB_LUT4 mux_56_Mux_0_i3_4_lut_4_lut (.I0(multi_byte_spi_trans_flag_r), 
            .I1(state[0]), .I2(state[1]), .I3(n19), .O(n3_adj_1373));
    defparam mux_56_Mux_0_i3_4_lut_4_lut.LUT_INIT = 16'hc131;
    SB_DFFE tx_shift_reg_i0_i15 (.Q(SDAT_c_15), .C(SLM_CLK_c), .E(n5081), 
            .D(n2330[15]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i43_4_lut_4_lut (.I0(state[2]), .I1(state[3]), .I2(state[1]), 
            .I3(state[0]), .O(n21));   // src/spi.v(88[9] 219[16])
    defparam i43_4_lut_4_lut.LUT_INIT = 16'hf01c;
    SB_LUT4 i3989_3_lut_4_lut (.I0(state[2]), .I1(state[3]), .I2(state[0]), 
            .I3(n3_adj_1373), .O(state_3__N_1122[0]));   // src/spi.v(88[9] 219[16])
    defparam i3989_3_lut_4_lut.LUT_INIT = 16'h1f0e;
    SB_DFF rx_shift_reg_i1 (.Q(\rx_shift_reg[1] ), .C(SLM_CLK_c), .D(n5706));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i2 (.Q(\rx_shift_reg[2] ), .C(SLM_CLK_c), .D(n5705));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i3 (.Q(\rx_shift_reg[3] ), .C(SLM_CLK_c), .D(n5704));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i4 (.Q(\rx_shift_reg[4] ), .C(SLM_CLK_c), .D(n5703));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i5 (.Q(\rx_shift_reg[5] ), .C(SLM_CLK_c), .D(n5702));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i6 (.Q(\rx_shift_reg[6] ), .C(SLM_CLK_c), .D(n5701));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i7 (.Q(\rx_shift_reg[7] ), .C(SLM_CLK_c), .D(n5700));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i1 (.Q(rx_buf_byte[1]), .C(SLM_CLK_c), .D(n5699));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i2 (.Q(rx_buf_byte[2]), .C(SLM_CLK_c), .D(n5698));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i3 (.Q(rx_buf_byte[3]), .C(SLM_CLK_c), .D(n5697));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i4 (.Q(rx_buf_byte[4]), .C(SLM_CLK_c), .D(n5696));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i5 (.Q(rx_buf_byte[5]), .C(SLM_CLK_c), .D(n5695));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i6 (.Q(rx_buf_byte[6]), .C(SLM_CLK_c), .D(n5694));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_1117_i2_3_lut (.I0(\tx_data_byte[1] ), .I1(\tx_shift_reg[0] ), 
            .I2(n2329), .I3(GND_net), .O(n2330[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_1117_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1117_i3_3_lut (.I0(\tx_data_byte[2] ), .I1(tx_shift_reg[1]), 
            .I2(n2329), .I3(GND_net), .O(n2330[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_1117_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1117_i4_3_lut (.I0(\tx_data_byte[3] ), .I1(tx_shift_reg[2]), 
            .I2(n2329), .I3(GND_net), .O(n2330[3]));   // src/spi.v(88[9] 219[16])
    defparam mux_1117_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1117_i5_3_lut (.I0(\tx_data_byte[4] ), .I1(tx_shift_reg[3]), 
            .I2(n2329), .I3(GND_net), .O(n2330[4]));   // src/spi.v(88[9] 219[16])
    defparam mux_1117_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF Rx_Recv_Byte_i7 (.Q(rx_buf_byte[7]), .C(SLM_CLK_c), .D(n5693));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_1117_i6_3_lut (.I0(\tx_data_byte[5] ), .I1(tx_shift_reg[4]), 
            .I2(n2329), .I3(GND_net), .O(n2330[5]));   // src/spi.v(88[9] 219[16])
    defparam mux_1117_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1117_i7_3_lut (.I0(\tx_data_byte[6] ), .I1(tx_shift_reg[5]), 
            .I2(n2329), .I3(GND_net), .O(n2330[6]));   // src/spi.v(88[9] 219[16])
    defparam mux_1117_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1117_i8_3_lut (.I0(\tx_data_byte[7] ), .I1(tx_shift_reg[6]), 
            .I2(n2329), .I3(GND_net), .O(n2330[7]));   // src/spi.v(88[9] 219[16])
    defparam mux_1117_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1117_i9_3_lut (.I0(tx_addr_byte[0]), .I1(tx_shift_reg[7]), 
            .I2(n2329), .I3(GND_net), .O(n2330[8]));   // src/spi.v(88[9] 219[16])
    defparam mux_1117_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1117_i10_3_lut (.I0(tx_addr_byte[1]), .I1(tx_shift_reg[8]), 
            .I2(n2329), .I3(GND_net), .O(n2330[9]));   // src/spi.v(88[9] 219[16])
    defparam mux_1117_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1139_9_lut (.I0(GND_net), .I1(multi_byte_counter[7]), .I2(n2406[6]), 
            .I3(n10312), .O(n315[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1139_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1117_i11_3_lut (.I0(tx_addr_byte[2]), .I1(tx_shift_reg[9]), 
            .I2(n2329), .I3(GND_net), .O(n2330[10]));   // src/spi.v(88[9] 219[16])
    defparam mux_1117_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1117_i12_3_lut (.I0(tx_addr_byte[3]), .I1(tx_shift_reg[10]), 
            .I2(n2329), .I3(GND_net), .O(n2330[11]));   // src/spi.v(88[9] 219[16])
    defparam mux_1117_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1117_i13_3_lut (.I0(tx_addr_byte[4]), .I1(tx_shift_reg[11]), 
            .I2(n2329), .I3(GND_net), .O(n2330[12]));   // src/spi.v(88[9] 219[16])
    defparam mux_1117_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1117_i14_3_lut (.I0(tx_addr_byte[5]), .I1(tx_shift_reg[12]), 
            .I2(n2329), .I3(GND_net), .O(n2330[13]));   // src/spi.v(88[9] 219[16])
    defparam mux_1117_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1117_i15_3_lut (.I0(tx_addr_byte[6]), .I1(tx_shift_reg[13]), 
            .I2(n2329), .I3(GND_net), .O(n2330[14]));   // src/spi.v(88[9] 219[16])
    defparam mux_1117_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF byte_recv_92_i3 (.Q(spi_rx_byte_ready), .C(SLM_CLK_c), .D(n1105[2]));   // src/spi.v(88[9] 219[16])
    SB_DFF byte_recv_92_i1 (.Q(SCK_c_0), .C(SLM_CLK_c), .D(n1105[0]));   // src/spi.v(88[9] 219[16])
    SB_LUT4 add_1139_8_lut (.I0(GND_net), .I1(multi_byte_counter[6]), .I2(n2406[6]), 
            .I3(n10311), .O(n315[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1139_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1139_8 (.CI(n10311), .I0(multi_byte_counter[6]), .I1(n2406[6]), 
            .CO(n10312));
    SB_LUT4 add_1139_7_lut (.I0(GND_net), .I1(multi_byte_counter[5]), .I2(n2406[6]), 
            .I3(n10310), .O(n315[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1139_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1139_7 (.CI(n10310), .I0(multi_byte_counter[5]), .I1(n2406[6]), 
            .CO(n10311));
    SB_LUT4 i4063_2_lut (.I0(n5199), .I1(state[3]), .I2(GND_net), .I3(GND_net), 
            .O(n5517));   // src/spi.v(76[8] 221[4])
    defparam i4063_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_72 (.I0(state[1]), .I1(n11370), .I2(n5009), .I3(state[3]), 
            .O(n5199));
    defparam i1_4_lut_adj_72.LUT_INIT = 16'h0a88;
    SB_LUT4 add_1139_6_lut (.I0(GND_net), .I1(multi_byte_counter[4]), .I2(n2406[6]), 
            .I3(n10309), .O(n315[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1139_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFE state_i3 (.Q(state[3]), .C(SLM_CLK_c), .E(n19_adj_1374), .D(state_3__N_1122[3]));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i2 (.Q(state[2]), .C(SLM_CLK_c), .E(n11091), .D(state_3__N_1122[2]));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i1 (.Q(state[1]), .C(SLM_CLK_c), .E(n5179), .D(state_3__N_1122[1]));   // src/spi.v(76[8] 221[4])
    SB_CARRY add_1139_6 (.CI(n10309), .I0(multi_byte_counter[4]), .I1(n2406[6]), 
            .CO(n10310));
    SB_LUT4 add_1139_5_lut (.I0(GND_net), .I1(multi_byte_counter[3]), .I2(n2406[6]), 
            .I3(n10308), .O(n315[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1139_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1139_5 (.CI(n10308), .I0(multi_byte_counter[3]), .I1(n2406[6]), 
            .CO(n10309));
    SB_DFFESR multi_byte_counter_i1 (.Q(multi_byte_counter[1]), .C(SLM_CLK_c), 
            .E(n5199), .D(n315[1]), .R(n5517));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i2 (.Q(multi_byte_counter[2]), .C(SLM_CLK_c), 
            .E(n5199), .D(n315[2]), .R(n5517));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i3 (.Q(multi_byte_counter[3]), .C(SLM_CLK_c), 
            .E(n5199), .D(n315[3]), .R(n5517));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i14 (.Q(tx_shift_reg[14]), .C(SLM_CLK_c), .E(n5081), 
            .D(n2330[14]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i13 (.Q(tx_shift_reg[13]), .C(SLM_CLK_c), .E(n5081), 
            .D(n2330[13]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i12 (.Q(tx_shift_reg[12]), .C(SLM_CLK_c), .E(n5081), 
            .D(n2330[12]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i11 (.Q(tx_shift_reg[11]), .C(SLM_CLK_c), .E(n5081), 
            .D(n2330[11]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i10 (.Q(tx_shift_reg[10]), .C(SLM_CLK_c), .E(n5081), 
            .D(n2330[10]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i9 (.Q(tx_shift_reg[9]), .C(SLM_CLK_c), .E(n5081), 
            .D(n2330[9]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i8 (.Q(tx_shift_reg[8]), .C(SLM_CLK_c), .E(n5081), 
            .D(n2330[8]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i7 (.Q(tx_shift_reg[7]), .C(SLM_CLK_c), .E(n5081), 
            .D(n2330[7]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i6 (.Q(tx_shift_reg[6]), .C(SLM_CLK_c), .E(n5081), 
            .D(n2330[6]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i5 (.Q(tx_shift_reg[5]), .C(SLM_CLK_c), .E(n5081), 
            .D(n2330[5]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i3_4_lut (.I0(state[3]), .I1(n5171), .I2(n11277), .I3(n5172), 
            .O(n5179));
    defparam i3_4_lut.LUT_INIT = 16'h4c00;
    SB_LUT4 i9907_2_lut (.I0(n19), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n11416));   // src/spi.v(88[9] 219[16])
    defparam i9907_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFE tx_shift_reg_i0_i4 (.Q(tx_shift_reg[4]), .C(SLM_CLK_c), .E(n5081), 
            .D(n2330[4]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i3 (.Q(tx_shift_reg[3]), .C(SLM_CLK_c), .E(n5081), 
            .D(n2330[3]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i2_3_lut (.I0(state[3]), .I1(n19), .I2(state[1]), .I3(GND_net), 
            .O(n11030));
    defparam i2_3_lut.LUT_INIT = 16'hbfbf;
    SB_DFFE tx_shift_reg_i0_i2 (.Q(tx_shift_reg[2]), .C(SLM_CLK_c), .E(n5081), 
            .D(n2330[2]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i1 (.Q(tx_shift_reg[1]), .C(SLM_CLK_c), .E(n5081), 
            .D(n2330[1]));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i4 (.Q(multi_byte_counter[4]), .C(SLM_CLK_c), 
            .E(n5199), .D(n315[4]), .R(n5517));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_56_Mux_1_i7_4_lut (.I0(n3), .I1(n11416), .I2(state[2]), 
            .I3(state[1]), .O(n7));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_1_i7_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 mux_56_Mux_1_i15_4_lut (.I0(n7), .I1(state[1]), .I2(state[3]), 
            .I3(state[0]), .O(state_3__N_1122[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_1_i15_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut (.I0(n5171), .I1(n11089), .I2(GND_net), .I3(GND_net), 
            .O(n11091));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_56_Mux_2_i3_3_lut (.I0(multi_byte_spi_trans_flag_r), .I1(state[0]), 
            .I2(state[1]), .I3(GND_net), .O(n3_adj_1375));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_2_i3_3_lut.LUT_INIT = 16'hc2c2;
    SB_LUT4 i4_4_lut (.I0(n11237), .I1(state[3]), .I2(spi_start_transfer_r), 
            .I3(state[0]), .O(n5172));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9660_2_lut (.I0(state[1]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n11237));
    defparam i9660_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESS multi_byte_counter_i5 (.Q(multi_byte_counter[5]), .C(SLM_CLK_c), 
            .E(n5199), .D(n315[5]), .S(n5517));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_56_Mux_2_i15_4_lut (.I0(n3_adj_1375), .I1(state[2]), .I2(state[3]), 
            .I3(state[0]), .O(state_3__N_1122[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_2_i15_4_lut.LUT_INIT = 16'hc2ce;
    SB_LUT4 i1_2_lut_adj_73 (.I0(n19), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_1376));
    defparam i1_2_lut_adj_73.LUT_INIT = 16'hdddd;
    SB_DFFESR multi_byte_counter_i6 (.Q(multi_byte_counter[6]), .C(SLM_CLK_c), 
            .E(n5199), .D(n315[6]), .R(n5517));   // src/spi.v(76[8] 221[4])
    SB_DFFESS multi_byte_counter_i7 (.Q(multi_byte_counter[7]), .C(SLM_CLK_c), 
            .E(n5199), .D(n315[7]), .S(n5517));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i1_4_lut_adj_74 (.I0(state[3]), .I1(n11089), .I2(n11237), 
            .I3(n4_adj_1376), .O(n11090));
    defparam i1_4_lut_adj_74.LUT_INIT = 16'h4c44;
    SB_LUT4 i3_4_lut_adj_75 (.I0(counter[0]), .I1(counter[1]), .I2(counter[2]), 
            .I3(counter[3]), .O(n11039));
    defparam i3_4_lut_adj_75.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_76 (.I0(n19), .I1(n21), .I2(GND_net), .I3(GND_net), 
            .O(n22));
    defparam i1_2_lut_adj_76.LUT_INIT = 16'h8888;
    SB_LUT4 i9956_4_lut (.I0(n22), .I1(n11273), .I2(n11277), .I3(state[3]), 
            .O(n19_adj_1374));
    defparam i9956_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 mux_56_Mux_3_i15_4_lut (.I0(n11418), .I1(state[1]), .I2(state[3]), 
            .I3(n2406[6]), .O(state_3__N_1122[3]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_3_i15_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i9997_3_lut (.I0(counter[4]), .I1(n11039), .I2(n4813), .I3(GND_net), 
            .O(n5113));   // src/spi.v(88[9] 219[16])
    defparam i9997_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_4_lut_4_lut (.I0(state[1]), .I1(state[3]), .I2(state[0]), 
            .I3(state[2]), .O(n5120));   // src/spi.v(88[9] 219[16])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h0140;
    SB_DFFE tx_shift_reg_i0_i0 (.Q(\tx_shift_reg[0] ), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n10792));   // src/spi.v(76[8] 221[4])
    SB_LUT4 add_1139_4_lut (.I0(GND_net), .I1(multi_byte_counter[2]), .I2(n2406[6]), 
            .I3(n10307), .O(n315[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1139_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1139_4 (.CI(n10307), .I0(multi_byte_counter[2]), .I1(n2406[6]), 
            .CO(n10308));
    SB_DFFESR counter_1347__i1 (.Q(counter[1]), .C(SLM_CLK_c), .E(n5142), 
            .D(n45[1]), .R(n5487));   // src/spi.v(183[28:41])
    SB_LUT4 i9901_3_lut (.I0(n2406[6]), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n11366));   // src/spi.v(88[9] 219[16])
    defparam i9901_3_lut.LUT_INIT = 16'hc4c4;
    SB_LUT4 mux_376_Mux_1_i7_4_lut (.I0(state[0]), .I1(state[2]), .I2(n19), 
            .I3(state[1]), .O(n7_adj_1377));   // src/spi.v(88[9] 219[16])
    defparam mux_376_Mux_1_i7_4_lut.LUT_INIT = 16'h02dd;
    SB_LUT4 mux_376_Mux_1_i15_4_lut (.I0(n7_adj_1377), .I1(n11366), .I2(state[3]), 
            .I3(state[2]), .O(n1105[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_376_Mux_1_i15_4_lut.LUT_INIT = 16'hfaca;
    SB_DFFESR counter_1347__i2 (.Q(counter[2]), .C(SLM_CLK_c), .E(n5142), 
            .D(n45[2]), .R(n5487));   // src/spi.v(183[28:41])
    SB_LUT4 add_1139_3_lut (.I0(GND_net), .I1(multi_byte_counter[1]), .I2(n2406[6]), 
            .I3(n10306), .O(n315[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1139_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR counter_1347__i3 (.Q(counter[3]), .C(SLM_CLK_c), .E(n5142), 
            .D(n45[3]), .R(n5487));   // src/spi.v(183[28:41])
    SB_CARRY add_1139_3 (.CI(n10306), .I0(multi_byte_counter[1]), .I1(n2406[6]), 
            .CO(n10307));
    SB_DFFESR counter_1347__i4 (.Q(counter[4]), .C(SLM_CLK_c), .E(n5142), 
            .D(n45[4]), .R(n5487));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1347__i5 (.Q(counter[5]), .C(SLM_CLK_c), .E(n5142), 
            .D(n45[5]), .R(n5487));   // src/spi.v(183[28:41])
    SB_LUT4 add_1139_2_lut (.I0(GND_net), .I1(multi_byte_counter[0]), .I2(n2406[6]), 
            .I3(GND_net), .O(n315[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1139_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_376_Mux_2_i15_4_lut_4_lut (.I0(state[0]), .I1(state[2]), 
            .I2(state[3]), .I3(state[1]), .O(n1105[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_376_Mux_2_i15_4_lut_4_lut.LUT_INIT = 16'h1008;
    SB_CARRY add_1139_2 (.CI(GND_net), .I0(multi_byte_counter[0]), .I1(n2406[6]), 
            .CO(n10306));
    SB_DFFESR counter_1347__i6 (.Q(counter[6]), .C(SLM_CLK_c), .E(n5142), 
            .D(n45[6]), .R(n5487));   // src/spi.v(183[28:41])
    SB_LUT4 i1_2_lut_4_lut (.I0(counter[0]), .I1(counter[1]), .I2(counter[3]), 
            .I3(counter[2]), .O(n8));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR counter_1347__i7 (.Q(counter[7]), .C(SLM_CLK_c), .E(n5142), 
            .D(n45[7]), .R(n5487));   // src/spi.v(183[28:41])
    SB_DFFESS counter_1347__i8 (.Q(counter[8]), .C(SLM_CLK_c), .E(n5142), 
            .D(n45[8]), .S(n5487));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1347__i9 (.Q(counter[9]), .C(SLM_CLK_c), .E(n5142), 
            .D(n45[9]), .R(n5487));   // src/spi.v(183[28:41])
    SB_DFF Rx_Recv_Byte_i0 (.Q(rx_buf_byte[0]), .C(SLM_CLK_c), .D(n5621));   // src/spi.v(76[8] 221[4])
    SB_LUT4 counter_1347_add_4_11_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[9]), 
            .I3(n10331), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1347_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1347_add_4_10_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[8]), 
            .I3(n10330), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1347_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1347_add_4_10 (.CI(n10330), .I0(VCC_net), .I1(counter[8]), 
            .CO(n10331));
    SB_LUT4 counter_1347_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[7]), 
            .I3(n10329), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1347_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1347_add_4_9 (.CI(n10329), .I0(VCC_net), .I1(counter[7]), 
            .CO(n10330));
    SB_LUT4 i9695_3_lut_4_lut (.I0(state[0]), .I1(state[2]), .I2(spi_start_transfer_r), 
            .I3(state[1]), .O(n11273));
    defparam i9695_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_77 (.I0(state[2]), .I1(state[3]), .I2(n19), 
            .I3(state[1]), .O(n5171));
    defparam i1_2_lut_4_lut_adj_77.LUT_INIT = 16'hefff;
    SB_DFFESR multi_byte_counter_i0 (.Q(multi_byte_counter[0]), .C(SLM_CLK_c), 
            .E(n5199), .D(n315[0]), .R(n5517));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i9883_4_lut (.I0(n8), .I1(state[1]), .I2(state[0]), .I3(state[2]), 
            .O(n11397));   // src/spi.v(88[9] 219[16])
    defparam i9883_4_lut.LUT_INIT = 16'hc08c;
    SB_LUT4 i1_4_lut_adj_78 (.I0(counter[4]), .I1(n11397), .I2(n11398), 
            .I3(state[3]), .O(n1105[0]));   // src/spi.v(88[9] 219[16])
    defparam i1_4_lut_adj_78.LUT_INIT = 16'ha088;
    SB_LUT4 i7_4_lut (.I0(multi_byte_counter[0]), .I1(n14_adj_1378), .I2(n10), 
            .I3(multi_byte_counter[6]), .O(n2406[6]));   // src/spi.v(208[21:52])
    defparam i7_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i9888_2_lut_3_lut (.I0(n19), .I1(state[0]), .I2(state[2]), 
            .I3(GND_net), .O(n11370));
    defparam i9888_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i10000_3_lut_4_lut (.I0(state[2]), .I1(state[0]), .I2(n24), 
            .I3(n16), .O(n5081));   // src/spi.v(88[9] 219[16])
    defparam i10000_3_lut_4_lut.LUT_INIT = 16'h000d;
    SB_LUT4 i3358_4_lut_4_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(state[3]), .O(n4813));   // src/spi.v(88[9] 219[16])
    defparam i3358_4_lut_4_lut_4_lut.LUT_INIT = 16'hfe75;
    SB_LUT4 i1_3_lut_4_lut (.I0(n2406[6]), .I1(state[0]), .I2(state[2]), 
            .I3(state[1]), .O(n5012));   // src/spi.v(88[9] 219[16])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i9887_2_lut_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(n8), .O(n11398));   // src/spi.v(88[9] 219[16])
    defparam i9887_2_lut_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i9670_2_lut (.I0(state[3]), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n11247));
    defparam i9670_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_79 (.I0(counter[1]), .I1(counter[3]), .I2(counter[2]), 
            .I3(GND_net), .O(n4931));
    defparam i2_3_lut_adj_79.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_2_lut (.I0(counter[7]), .I1(counter[5]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_1379));   // src/spi.v(141[21:41])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(counter[4]), .I1(counter[6]), .I2(counter[8]), 
            .I3(counter[9]), .O(n14_adj_1380));   // src/spi.v(141[21:41])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_80 (.I0(counter[0]), .I1(n14_adj_1380), .I2(n10_adj_1379), 
            .I3(n4931), .O(n19));   // src/spi.v(141[21:41])
    defparam i7_4_lut_adj_80.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_adj_81 (.I0(state[0]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5009));   // src/spi.v(88[9] 219[16])
    defparam i1_2_lut_adj_81.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_82 (.I0(multi_byte_counter[2]), .I1(multi_byte_counter[4]), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // src/spi.v(208[21:52])
    defparam i2_2_lut_adj_82.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_83 (.I0(multi_byte_counter[3]), .I1(multi_byte_counter[1]), 
            .I2(multi_byte_counter[5]), .I3(multi_byte_counter[7]), .O(n14_adj_1378));   // src/spi.v(208[21:52])
    defparam i6_4_lut_adj_83.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut (.I0(state[3]), .I1(state[0]), .I2(state[2]), 
            .I3(GND_net), .O(n14));   // src/spi.v(88[9] 219[16])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf1f1;
    SB_LUT4 i1_3_lut_4_lut_adj_84 (.I0(state[0]), .I1(state[2]), .I2(n11030), 
            .I3(n5172), .O(n11089));
    defparam i1_3_lut_4_lut_adj_84.LUT_INIT = 16'hf700;
    
endmodule
//
// Verilog Description of module usb3_if
//

module usb3_if (reset_per_frame, SLM_CLK_c, DEBUG_9_c, VCC_net, FT_RD_c, 
            FIFO_CLK_c, DEBUG_3_c_0, dc32_fifo_write_enable, buffer_switch_done, 
            buffer_switch_done_latched, FT_OE_c, FR_RXF_c, GND_net, 
            DEBUG_1_c, FIFO_D0_c_0) /* synthesis syn_module_defined=1 */ ;
    input reset_per_frame;
    input SLM_CLK_c;
    input DEBUG_9_c;
    input VCC_net;
    output FT_RD_c;
    input FIFO_CLK_c;
    output DEBUG_3_c_0;
    output dc32_fifo_write_enable;
    input buffer_switch_done;
    output buffer_switch_done_latched;
    output FT_OE_c;
    input FR_RXF_c;
    input GND_net;
    input DEBUG_1_c;
    input FIFO_D0_c_0;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    
    wire reset_per_frame_latched, dc32_fifo_empty_latched, FT_RD_N_500, 
        n2603, n5069;
    wire [4:0]state_timeout_counter;   // src/usb3_if.v(64[11:32])
    
    wire n9407;
    wire [6:0]n70;
    
    wire n5278;
    wire [5:0]num_words_curr_line;   // src/usb3_if.v(60[11:30])
    
    wire n9417;
    wire [31:0]dc32_fifo_data_in_latched;   // src/usb3_if.v(66[12:37])
    
    wire write_to_dc32_fifo_latched;
    wire [5:0]num_words_curr_line_5__N_434;
    
    wire FT_OE_N_489, n2604, n8065;
    wire [15:0]n650;
    
<<<<<<< HEAD
    wire FT_OE_N_495, write_to_dc32_fifo_latched_N_502, n2605, n2606;
    wire [10:0]num_lines_clocked_out_10__N_440;
    
    wire n5254;
    wire [10:0]num_lines_clocked_out;   // src/usb3_if.v(63[12:33])
    
    wire n3410;
    wire [3:0]n154;
    
    wire n607, n2623, n63, n10290, n71, n10230, n10228, n10231, 
        n10232, n10229, n10289, n709, n64, n10288, n10237, n10287, 
        n10286, n10236, n10235, n10234, n706, n10233, n3378, n3385, 
        n696, n3390, n11042, n9411, n139, n5660, n2617, n2620, 
        n8, n609, FT_OE_N_494, n11384, n10424, n6, n2609, n18, 
        n16, n20, n4644, FT_OE_N_490, n73_adj_1369, n3391, n605, 
        n623, n4997, n2602, n11139, n10978, n16_adj_1370, n69, 
        n6_adj_1371, n11701, n4270, n11051, n7, n85, n6_adj_1372, 
        n10;
    
    SB_DFF reset_per_frame_latched_108 (.Q(reset_per_frame_latched), .C(SLM_CLK_c), 
           .D(reset_per_frame));   // src/usb3_if.v(70[8] 83[4])
    SB_DFF dc32_fifo_empty_latched_109 (.Q(dc32_fifo_empty_latched), .C(SLM_CLK_c), 
           .D(DEBUG_9_c));   // src/usb3_if.v(70[8] 83[4])
    SB_DFFESS FT_RD_111 (.Q(FT_RD_c), .C(FIFO_CLK_c), .E(VCC_net), .D(FT_RD_N_500), 
            .S(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(FIFO_CLK_c), 
            .E(n5069), .D(n2603), .R(n9407));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_words_curr_line_i1 (.Q(num_words_curr_line[1]), .C(FIFO_CLK_c), 
            .E(n5278), .D(n70[1]), .R(n9417));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_words_curr_line_i2 (.Q(num_words_curr_line[2]), .C(FIFO_CLK_c), 
            .E(n5278), .D(n70[2]), .R(n9417));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFN dc32_fifo_data_in_i1 (.Q(DEBUG_3_c_0), .C(FIFO_CLK_c), .D(dc32_fifo_data_in_latched[0]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN write_to_dc32_fifo_119 (.Q(dc32_fifo_write_enable), .C(FIFO_CLK_c), 
            .D(write_to_dc32_fifo_latched));   // src/usb3_if.v(204[8] 207[4])
    SB_DFF buffer_switch_done_latched_107 (.Q(buffer_switch_done_latched), 
           .C(SLM_CLK_c), .D(buffer_switch_done));   // src/usb3_if.v(70[8] 83[4])
    SB_DFFESS num_words_curr_line_i3 (.Q(num_words_curr_line[3]), .C(FIFO_CLK_c), 
            .E(n5278), .D(num_words_curr_line_5__N_434[3]), .S(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESS FT_OE_110 (.Q(FT_OE_c), .C(FIFO_CLK_c), .E(VCC_net), .D(FT_OE_N_489), 
            .S(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESS state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(FIFO_CLK_c), 
            .E(n5069), .D(n2604), .S(n9407));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i244_4_lut (.I0(n8065), .I1(FR_RXF_c), .I2(n650[5]), .I3(FT_OE_N_495), 
            .O(write_to_dc32_fifo_latched_N_502));   // src/usb3_if.v(97[9] 199[16])
    defparam i244_4_lut.LUT_INIT = 16'h3a0a;
    SB_DFFESR state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(FIFO_CLK_c), 
            .E(n5069), .D(n2605), .R(n9407));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_words_curr_line_i4 (.Q(num_words_curr_line[4]), .C(FIFO_CLK_c), 
            .E(n5278), .D(n70[4]), .R(n9417));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(FIFO_CLK_c), 
            .E(n5069), .D(n2606), .R(n9407));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESS num_words_curr_line_i5 (.Q(num_words_curr_line[5]), .C(FIFO_CLK_c), 
            .E(n5278), .D(num_words_curr_line_5__N_434[5]), .S(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i1 (.Q(num_lines_clocked_out[1]), .C(FIFO_CLK_c), 
            .E(n5254), .D(num_lines_clocked_out_10__N_440[1]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i2 (.Q(num_lines_clocked_out[2]), .C(FIFO_CLK_c), 
            .E(n5254), .D(num_lines_clocked_out_10__N_440[2]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFSS state_FSM_i1 (.Q(n650[0]), .C(FIFO_CLK_c), .D(n3410), .S(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFESR num_lines_clocked_out_i3 (.Q(num_lines_clocked_out[3]), .C(FIFO_CLK_c), 
            .E(n5254), .D(num_lines_clocked_out_10__N_440[3]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i4 (.Q(num_lines_clocked_out[4]), .C(FIFO_CLK_c), 
            .E(n5254), .D(num_lines_clocked_out_10__N_440[4]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i5 (.Q(num_lines_clocked_out[5]), .C(FIFO_CLK_c), 
            .E(n5254), .D(num_lines_clocked_out_10__N_440[5]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i6 (.Q(num_lines_clocked_out[6]), .C(FIFO_CLK_c), 
            .E(n5254), .D(num_lines_clocked_out_10__N_440[6]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFSR write_to_dc32_fifo_latched_113 (.Q(write_to_dc32_fifo_latched), 
            .C(FIFO_CLK_c), .D(write_to_dc32_fifo_latched_N_502), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESS num_lines_clocked_out_i7 (.Q(num_lines_clocked_out[7]), .C(FIFO_CLK_c), 
            .E(n5254), .D(num_lines_clocked_out_10__N_440[7]), .S(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i8 (.Q(num_lines_clocked_out[8]), .C(FIFO_CLK_c), 
            .E(n5254), .D(num_lines_clocked_out_10__N_440[8]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i9 (.Q(num_lines_clocked_out[9]), .C(FIFO_CLK_c), 
            .E(n5254), .D(num_lines_clocked_out_10__N_440[9]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i10 (.Q(num_lines_clocked_out[10]), .C(FIFO_CLK_c), 
            .E(n5254), .D(num_lines_clocked_out_10__N_440[10]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i1966_4_lut (.I0(n650[0]), .I1(n154[0]), .I2(n607), .I3(n2623), 
            .O(n3410));   // src/usb3_if.v(97[9] 199[16])
    defparam i1966_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 sub_114_add_2_7_lut (.I0(n71), .I1(num_words_curr_line[5]), 
            .I2(VCC_net), .I3(n10290), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_114_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_116_add_2_5_lut (.I0(GND_net), .I1(num_lines_clocked_out[3]), 
            .I2(VCC_net), .I3(n10230), .O(num_lines_clocked_out_10__N_440[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_116_add_2_3_lut (.I0(GND_net), .I1(num_lines_clocked_out[1]), 
            .I2(VCC_net), .I3(n10228), .O(num_lines_clocked_out_10__N_440[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_116_add_2_6 (.CI(n10231), .I0(num_lines_clocked_out[4]), 
            .I1(VCC_net), .CO(n10232));
    SB_CARRY sub_116_add_2_3 (.CI(n10228), .I0(num_lines_clocked_out[1]), 
            .I1(VCC_net), .CO(n10229));
    SB_LUT4 sub_114_add_2_6_lut (.I0(GND_net), .I1(num_words_curr_line[4]), 
            .I2(VCC_net), .I3(n10289), .O(n70[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_114_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_114_add_2_6 (.CI(n10289), .I0(num_words_curr_line[4]), 
            .I1(VCC_net), .CO(n10290));
    SB_LUT4 sub_116_add_2_7_lut (.I0(GND_net), .I1(num_lines_clocked_out[5]), 
            .I2(VCC_net), .I3(n10232), .O(num_lines_clocked_out_10__N_440[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR state_FSM_i9 (.Q(n650[8]), .C(FIFO_CLK_c), .D(n709), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_LUT4 sub_114_add_2_5_lut (.I0(n71), .I1(num_words_curr_line[3]), 
            .I2(VCC_net), .I3(n10288), .O(n64)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_114_add_2_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_116_add_2_12_lut (.I0(GND_net), .I1(num_lines_clocked_out[10]), 
            .I2(VCC_net), .I3(n10237), .O(num_lines_clocked_out_10__N_440[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_114_add_2_5 (.CI(n10288), .I0(num_words_curr_line[3]), 
            .I1(VCC_net), .CO(n10289));
    SB_CARRY sub_116_add_2_5 (.CI(n10230), .I0(num_lines_clocked_out[3]), 
            .I1(VCC_net), .CO(n10231));
    SB_LUT4 sub_114_add_2_4_lut (.I0(GND_net), .I1(num_words_curr_line[2]), 
            .I2(VCC_net), .I3(n10287), .O(n70[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_114_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_114_add_2_4 (.CI(n10287), .I0(num_words_curr_line[2]), 
            .I1(VCC_net), .CO(n10288));
    SB_LUT4 sub_114_add_2_3_lut (.I0(GND_net), .I1(num_words_curr_line[1]), 
            .I2(VCC_net), .I3(n10286), .O(n70[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_114_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_116_add_2_6_lut (.I0(GND_net), .I1(num_lines_clocked_out[4]), 
            .I2(VCC_net), .I3(n10231), .O(num_lines_clocked_out_10__N_440[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_116_add_2_11_lut (.I0(GND_net), .I1(num_lines_clocked_out[9]), 
            .I2(VCC_net), .I3(n10236), .O(num_lines_clocked_out_10__N_440[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_116_add_2_11 (.CI(n10236), .I0(num_lines_clocked_out[9]), 
            .I1(VCC_net), .CO(n10237));
    SB_LUT4 sub_116_add_2_10_lut (.I0(GND_net), .I1(num_lines_clocked_out[8]), 
            .I2(VCC_net), .I3(n10235), .O(num_lines_clocked_out_10__N_440[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_116_add_2_10 (.CI(n10235), .I0(num_lines_clocked_out[8]), 
            .I1(VCC_net), .CO(n10236));
    SB_CARRY sub_114_add_2_3 (.CI(n10286), .I0(num_words_curr_line[1]), 
            .I1(VCC_net), .CO(n10287));
    SB_LUT4 sub_114_add_2_2_lut (.I0(GND_net), .I1(num_words_curr_line[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n70[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_114_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_114_add_2_2 (.CI(VCC_net), .I0(num_words_curr_line[0]), 
            .I1(GND_net), .CO(n10286));
    SB_LUT4 sub_116_add_2_9_lut (.I0(GND_net), .I1(num_lines_clocked_out[7]), 
            .I2(VCC_net), .I3(n10234), .O(num_lines_clocked_out_10__N_440[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR state_FSM_i8 (.Q(n650[7]), .C(FIFO_CLK_c), .D(n706), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_CARRY sub_116_add_2_7 (.CI(n10232), .I0(num_lines_clocked_out[5]), 
            .I1(VCC_net), .CO(n10233));
    SB_DFFSR state_FSM_i7 (.Q(n650[6]), .C(FIFO_CLK_c), .D(n3378), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFSR state_FSM_i6 (.Q(n650[5]), .C(FIFO_CLK_c), .D(n3385), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFSR state_FSM_i4 (.Q(n650[3]), .C(FIFO_CLK_c), .D(n696), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFSR state_FSM_i3 (.Q(n650[2]), .C(FIFO_CLK_c), .D(n3390), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFSR state_FSM_i2 (.Q(n650[1]), .C(FIFO_CLK_c), .D(n11042), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_CARRY sub_116_add_2_9 (.CI(n10234), .I0(num_lines_clocked_out[7]), 
            .I1(VCC_net), .CO(n10235));
    SB_LUT4 sub_116_add_2_8_lut (.I0(GND_net), .I1(num_lines_clocked_out[6]), 
            .I2(VCC_net), .I3(n10233), .O(num_lines_clocked_out_10__N_440[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut (.I0(n63), .I1(n9411), .I2(GND_net), .I3(GND_net), 
            .O(num_words_curr_line_5__N_434[5]));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY sub_116_add_2_8 (.CI(n10233), .I0(num_lines_clocked_out[6]), 
            .I1(VCC_net), .CO(n10234));
    SB_LUT4 sub_116_add_2_4_lut (.I0(GND_net), .I1(num_lines_clocked_out[2]), 
            .I2(VCC_net), .I3(n10229), .O(num_lines_clocked_out_10__N_440[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_116_add_2_2_lut (.I0(GND_net), .I1(num_lines_clocked_out[0]), 
            .I2(n139), .I3(VCC_net), .O(num_lines_clocked_out_10__N_440[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF state_FSM_i5 (.Q(n650[4]), .C(FIFO_CLK_c), .D(n5660));   // src/usb3_if.v(97[9] 199[16])
    SB_LUT4 i1_2_lut_adj_49 (.I0(reset_per_frame_latched), .I1(n650[3]), 
            .I2(GND_net), .I3(GND_net), .O(n5660));   // src/usb3_if.v(70[8] 83[4])
    defparam i1_2_lut_adj_49.LUT_INIT = 16'h4444;
    SB_LUT4 mux_1297_i5_4_lut (.I0(n2617), .I1(state_timeout_counter[4]), 
            .I2(n2620), .I3(n8), .O(n2606));   // src/usb3_if.v(97[9] 199[16])
    defparam mux_1297_i5_4_lut.LUT_INIT = 16'hca3a;
    SB_LUT4 i6457_2_lut (.I0(n154[0]), .I1(n2623), .I2(GND_net), .I3(GND_net), 
            .O(n2617));   // src/usb3_if.v(173[26] 175[24])
    defparam i6457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i9873_3_lut_4_lut (.I0(n609), .I1(n650[2]), .I2(n139), .I3(FT_OE_N_494), 
            .O(n11384));   // src/usb3_if.v(97[9] 199[16])
    defparam i9873_3_lut_4_lut.LUT_INIT = 16'h4404;
    SB_LUT4 i2_3_lut_4_lut (.I0(n650[0]), .I1(n650[2]), .I2(n650[6]), 
            .I3(n650[1]), .O(n10424));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1297_i4_4_lut (.I0(n2617), .I1(state_timeout_counter[3]), 
            .I2(n2620), .I3(n6), .O(n2605));   // src/usb3_if.v(97[9] 199[16])
    defparam mux_1297_i4_4_lut.LUT_INIT = 16'hca3a;
    SB_LUT4 i1842_3_lut_3_lut (.I0(n650[0]), .I1(n650[2]), .I2(n650[5]), 
            .I3(GND_net), .O(n2609));
    defparam i1842_3_lut_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 i1_2_lut_3_lut (.I0(n650[5]), .I1(FT_OE_N_495), .I2(DEBUG_1_c), 
            .I3(GND_net), .O(n71));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i7_4_lut (.I0(num_lines_clocked_out[7]), .I1(num_lines_clocked_out[2]), 
            .I2(num_lines_clocked_out[9]), .I3(num_lines_clocked_out[0]), 
            .O(n18));   // src/usb3_if.v(164[29:57])
    defparam i7_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i5_2_lut (.I0(num_lines_clocked_out[1]), .I1(num_lines_clocked_out[5]), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // src/usb3_if.v(164[29:57])
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut (.I0(num_lines_clocked_out[6]), .I1(n18), .I2(num_lines_clocked_out[3]), 
            .I3(num_lines_clocked_out[10]), .O(n20));   // src/usb3_if.v(164[29:57])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(num_lines_clocked_out[4]), .I1(n20), .I2(n16), 
            .I3(num_lines_clocked_out[8]), .O(n154[0]));   // src/usb3_if.v(164[29:57])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1297_i3_4_lut (.I0(n2623), .I1(n4644), .I2(n2620), .I3(n154[0]), 
            .O(n2604));   // src/usb3_if.v(97[9] 199[16])
    defparam mux_1297_i3_4_lut.LUT_INIT = 16'h3f35;
    SB_LUT4 i259_4_lut (.I0(FT_OE_N_490), .I1(n8065), .I2(n10424), .I3(n650[5]), 
            .O(FT_OE_N_489));   // src/usb3_if.v(97[9] 199[16])
    defparam i259_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i1_4_lut (.I0(n650[5]), .I1(FT_OE_N_494), .I2(n650[3]), .I3(n139), 
            .O(n9411));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_4_lut.LUT_INIT = 16'h5051;
    SB_LUT4 i1_2_lut_adj_50 (.I0(n64), .I1(n9411), .I2(GND_net), .I3(GND_net), 
            .O(num_words_curr_line_5__N_434[3]));
    defparam i1_2_lut_adj_50.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_51 (.I0(n73_adj_1369), .I1(n650[1]), .I2(GND_net), 
            .I3(GND_net), .O(n3391));   // src/usb3_if.v(153[17] 176[20])
    defparam i1_2_lut_adj_51.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_52 (.I0(n2617), .I1(n605), .I2(n3391), .I3(n650[0]), 
            .O(n11042));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_4_lut_adj_52.LUT_INIT = 16'hfefa;
    SB_LUT4 i1947_4_lut (.I0(n650[2]), .I1(FT_OE_N_495), .I2(n623), .I3(n650[5]), 
            .O(n3390));   // src/usb3_if.v(97[9] 199[16])
    defparam i1947_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 i1_2_lut_adj_53 (.I0(n650[1]), .I1(n73_adj_1369), .I2(GND_net), 
            .I3(GND_net), .O(n696));   // src/usb3_if.v(153[21:49])
    defparam i1_2_lut_adj_53.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_54 (.I0(n650[5]), .I1(FT_OE_N_495), .I2(GND_net), 
            .I3(GND_net), .O(n4997));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_2_lut_adj_54.LUT_INIT = 16'h8888;
    SB_LUT4 i173_3_lut_3_lut_4_lut (.I0(FT_OE_N_495), .I1(DEBUG_1_c), .I2(n609), 
            .I3(DEBUG_9_c), .O(n623));   // src/usb3_if.v(153[17] 176[20])
    defparam i173_3_lut_3_lut_4_lut.LUT_INIT = 16'hf8fd;
    SB_CARRY sub_116_add_2_2 (.CI(VCC_net), .I0(num_lines_clocked_out[0]), 
            .I1(n139), .CO(n10228));
    SB_LUT4 i1935_4_lut (.I0(n73_adj_1369), .I1(FR_RXF_c), .I2(n650[6]), 
            .I3(n4997), .O(n3378));   // src/usb3_if.v(97[9] 199[16])
    defparam i1935_4_lut.LUT_INIT = 16'heca0;
    SB_LUT4 mux_1297_i1_3_lut (.I0(n2623), .I1(state_timeout_counter[0]), 
            .I2(n2620), .I3(GND_net), .O(n2602));   // src/usb3_if.v(97[9] 199[16])
    defparam mux_1297_i1_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_3_lut (.I0(n609), .I1(FR_RXF_c), .I2(DEBUG_1_c), .I3(GND_net), 
            .O(n73_adj_1369));   // src/usb3_if.v(153[17] 176[20])
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_55 (.I0(n650[6]), .I1(n73_adj_1369), .I2(GND_net), 
            .I3(GND_net), .O(n706));   // src/usb3_if.v(153[21:49])
    defparam i1_2_lut_adj_55.LUT_INIT = 16'h2222;
    SB_LUT4 i157_2_lut_3_lut (.I0(buffer_switch_done_latched), .I1(dc32_fifo_empty_latched), 
            .I2(FR_RXF_c), .I3(GND_net), .O(n607));   // src/usb3_if.v(99[21:96])
    defparam i157_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i155_2_lut_3_lut (.I0(buffer_switch_done_latched), .I1(dc32_fifo_empty_latched), 
            .I2(FR_RXF_c), .I3(GND_net), .O(n605));   // src/usb3_if.v(99[21:96])
    defparam i155_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i9563_2_lut (.I0(n650[2]), .I1(n650[5]), .I2(GND_net), .I3(GND_net), 
            .O(n11139));
    defparam i9563_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_56 (.I0(reset_per_frame_latched), .I1(n650[4]), 
            .I2(n11139), .I3(n650[6]), .O(n10978));   // src/usb3_if.v(59[5:28])
    defparam i1_4_lut_adj_56.LUT_INIT = 16'haaab;
    SB_LUT4 i23_4_lut (.I0(n11384), .I1(FT_OE_N_490), .I2(n650[5]), .I3(n650[3]), 
            .O(n16_adj_1370));
    defparam i23_4_lut.LUT_INIT = 16'h3f3a;
    SB_LUT4 i1_2_lut_3_lut_adj_57 (.I0(FT_OE_N_495), .I1(DEBUG_1_c), .I2(n650[3]), 
            .I3(GND_net), .O(n69));   // src/usb3_if.v(154[25:87])
    defparam i1_2_lut_3_lut_adj_57.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_adj_58 (.I0(reset_per_frame_latched), .I1(n650[6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_1371));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_2_lut_adj_58.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_59 (.I0(n650[7]), .I1(n8065), .I2(GND_net), .I3(GND_net), 
            .O(n709));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_2_lut_adj_59.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(n650[5]), .I1(n650[4]), .I2(n650[2]), .I3(n6_adj_1371), 
            .O(n11701));   // src/usb3_if.v(97[9] 199[16])
    defparam i4_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i9621_4_lut (.I0(reset_per_frame_latched), .I1(n650[5]), .I2(n16_adj_1370), 
            .I3(n69), .O(n9417));   // src/usb3_if.v(59[5:28])
    defparam i9621_4_lut.LUT_INIT = 16'hbaaa;
    SB_LUT4 i1942_3_lut_4_lut (.I0(FR_RXF_c), .I1(n650[4]), .I2(n650[8]), 
            .I3(n4997), .O(n3385));   // src/usb3_if.v(97[9] 199[16])
    defparam i1942_3_lut_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i1_2_lut_adj_60 (.I0(reset_per_frame_latched), .I1(n16_adj_1370), 
            .I2(GND_net), .I3(GND_net), .O(n5278));
    defparam i1_2_lut_adj_60.LUT_INIT = 16'heeee;
    SB_CARRY sub_116_add_2_4 (.CI(n10229), .I0(num_lines_clocked_out[2]), 
            .I1(VCC_net), .CO(n10230));
    SB_LUT4 i1_3_lut_4_lut (.I0(FT_OE_N_494), .I1(n609), .I2(n650[2]), 
            .I3(reset_per_frame_latched), .O(n5254));   // src/usb3_if.v(153[17] 176[20])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hff10;
    SB_LUT4 i2_3_lut_4_lut_adj_61 (.I0(FT_OE_N_494), .I1(n609), .I2(n139), 
            .I3(n650[2]), .O(n2623));   // src/usb3_if.v(153[17] 176[20])
    defparam i2_3_lut_4_lut_adj_61.LUT_INIT = 16'h0100;
    SB_LUT4 i6619_2_lut_3_lut_4_lut (.I0(n609), .I1(n650[2]), .I2(FT_OE_N_495), 
            .I3(DEBUG_1_c), .O(n8065));   // src/usb3_if.v(97[9] 199[16])
    defparam i6619_2_lut_3_lut_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i1483_2_lut_4_lut (.I0(state_timeout_counter[3]), .I1(state_timeout_counter[1]), 
            .I2(state_timeout_counter[0]), .I3(state_timeout_counter[2]), 
            .O(n8));   // src/usb3_if.v(179[42:69])
    defparam i1483_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR dc32_fifo_data_in_latched__i0 (.Q(dc32_fifo_data_in_latched[0]), 
            .C(FIFO_CLK_c), .E(n11701), .D(FIFO_D0_c_0), .R(n10978));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i9949_2_lut (.I0(FT_OE_N_495), .I1(DEBUG_9_c), .I2(GND_net), 
            .I3(GND_net), .O(n139));   // src/usb3_if.v(161[30:87])
    defparam i9949_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1841_3_lut (.I0(FR_RXF_c), .I1(FT_OE_N_495), .I2(n650[2]), 
            .I3(GND_net), .O(n4270));   // src/usb3_if.v(97[9] 199[16])
    defparam i1841_3_lut.LUT_INIT = 16'hc5c5;
    SB_DFFESR num_lines_clocked_out_i0 (.Q(num_lines_clocked_out[0]), .C(FIFO_CLK_c), 
            .E(n5254), .D(num_lines_clocked_out_10__N_440[0]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i1962_3_lut (.I0(n609), .I1(DEBUG_1_c), .I2(n4270), .I3(GND_net), 
            .O(n2620));   // src/usb3_if.v(97[9] 199[16])
    defparam i1962_3_lut.LUT_INIT = 16'hbaba;
    SB_DFFESR num_words_curr_line_i0 (.Q(num_words_curr_line[0]), .C(FIFO_CLK_c), 
            .E(n5278), .D(n70[0]), .R(n9417));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(FIFO_CLK_c), 
            .E(n5069), .D(n2602), .R(n9407));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i1_4_lut_adj_62 (.I0(n650[5]), .I1(n650[0]), .I2(FT_OE_N_490), 
            .I3(n605), .O(n11051));   // src/usb3_if.v(154[25:87])
    defparam i1_4_lut_adj_62.LUT_INIT = 16'h0ace;
    SB_LUT4 i4_4_lut_adj_63 (.I0(n7), .I1(n11051), .I2(n650[3]), .I3(n650[7]), 
            .O(n85));   // src/usb3_if.v(154[25:87])
    defparam i4_4_lut_adj_63.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_64 (.I0(reset_per_frame_latched), .I1(n2609), .I2(n85), 
            .I3(GND_net), .O(n9407));   // src/usb3_if.v(70[8] 83[4])
    defparam i1_3_lut_adj_64.LUT_INIT = 16'h0404;
    SB_LUT4 i9967_2_lut (.I0(reset_per_frame_latched), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n5069));
    defparam i9967_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 mux_1297_i2_4_lut (.I0(n2623), .I1(state_timeout_counter[1]), 
            .I2(n2620), .I3(state_timeout_counter[0]), .O(n2603));   // src/usb3_if.v(97[9] 199[16])
    defparam mux_1297_i2_4_lut.LUT_INIT = 16'hca3a;
    SB_LUT4 i1_2_lut_adj_65 (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_1372));   // src/usb3_if.v(153[21:49])
    defparam i1_2_lut_adj_65.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_66 (.I0(state_timeout_counter[3]), .I1(state_timeout_counter[2]), 
            .I2(state_timeout_counter[0]), .I3(n6_adj_1372), .O(n609));   // src/usb3_if.v(153[21:49])
    defparam i4_4_lut_adj_66.LUT_INIT = 16'hffef;
    SB_LUT4 FT_OE_I_8_2_lut (.I0(FT_OE_N_495), .I1(DEBUG_1_c), .I2(GND_net), 
            .I3(GND_net), .O(FT_OE_N_494));   // src/usb3_if.v(154[25:87])
    defparam FT_OE_I_8_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut_adj_67 (.I0(num_words_curr_line[2]), .I1(num_words_curr_line[5]), 
            .I2(num_words_curr_line[0]), .I3(num_words_curr_line[1]), .O(n10));   // src/usb3_if.v(132[21:47])
    defparam i4_4_lut_adj_67.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(num_words_curr_line[3]), .I1(n10), .I2(num_words_curr_line[4]), 
            .I3(GND_net), .O(FT_OE_N_495));   // src/usb3_if.v(132[21:47])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_2_lut (.I0(n650[4]), .I1(n650[8]), .I2(GND_net), .I3(GND_net), 
            .O(n7));   // src/usb3_if.v(154[25:87])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6341_2_lut (.I0(FR_RXF_c), .I1(FT_OE_N_495), .I2(GND_net), 
            .I3(GND_net), .O(FT_OE_N_490));   // src/usb3_if.v(137[22] 148[20])
    defparam i6341_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1873_4_lut (.I0(n8065), .I1(FT_OE_N_490), .I2(n650[5]), .I3(n7), 
            .O(FT_RD_N_500));   // src/usb3_if.v(97[9] 199[16])
    defparam i1873_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 i1_2_lut_3_lut_adj_68 (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[0]), 
            .I2(state_timeout_counter[2]), .I3(GND_net), .O(n4644));   // src/usb3_if.v(179[42:69])
    defparam i1_2_lut_3_lut_adj_68.LUT_INIT = 16'h1e1e;
    SB_LUT4 i1475_2_lut_3_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[0]), 
            .I2(state_timeout_counter[2]), .I3(GND_net), .O(n6));   // src/usb3_if.v(179[42:69])
    defparam i1475_2_lut_3_lut.LUT_INIT = 16'hfefe;
=======
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10856 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_5 ), 
            .I2(\REG.mem_15_5 ), .I3(rd_addr_r_c[1]), .O(n12773));
    defparam rd_addr_r_0__bdd_4_lut_10856.LUT_INIT = 16'he4aa;
    SB_LUT4 n13421_bdd_4_lut (.I0(n13421), .I1(n11523), .I2(n11522), .I3(rd_addr_r_c[2]), 
            .O(n13424));
    defparam n13421_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4395_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_51_6 ), .O(n5778));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4395_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFSR \afull_flag_impl.af_flag_ext_r_121  (.Q(dc32_fifo_almost_full), 
            .C(FIFO_CLK_c), .D(\afull_flag_impl.af_flag_nxt_w ), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(410[29] 422[32])
    SB_LUT4 n12773_bdd_4_lut (.I0(n12773), .I1(\REG.mem_13_5 ), .I2(\REG.mem_12_5 ), 
            .I3(rd_addr_r_c[1]), .O(n12776));
    defparam n12773_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4394_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_51_5 ), .O(n5777));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4394_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4393_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_51_4 ), .O(n5776));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4393_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10851 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_0 ), 
            .I2(\REG.mem_31_0 ), .I3(rd_addr_r_c[1]), .O(n12767));
    defparam rd_addr_r_0__bdd_4_lut_10851.LUT_INIT = 16'he4aa;
    SB_LUT4 n12767_bdd_4_lut (.I0(n12767), .I1(\REG.mem_29_0 ), .I2(\REG.mem_28_0 ), 
            .I3(rd_addr_r_c[1]), .O(n12770));
    defparam n12767_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9184_3_lut (.I0(n13724), .I1(n13700), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11022));
    defparam i9184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4392_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_51_3 ), .O(n5775));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4392_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11405 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_13 ), 
            .I2(\REG.mem_55_13 ), .I3(rd_addr_r_c[1]), .O(n13415));
    defparam rd_addr_r_0__bdd_4_lut_11405.LUT_INIT = 16'he4aa;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i3_1_lut (.I0(rd_addr_r_c[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4094_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_34_2 ), .O(n5477));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4094_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9592_3_lut (.I0(\REG.mem_38_7 ), .I1(\REG.mem_39_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11430));
    defparam i9592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9591_3_lut (.I0(\REG.mem_36_7 ), .I1(\REG.mem_37_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11429));
    defparam i9591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9555_3_lut (.I0(\REG.mem_16_8 ), .I1(\REG.mem_17_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11393));
    defparam i9555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9556_3_lut (.I0(\REG.mem_18_8 ), .I1(\REG.mem_19_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11394));
    defparam i9556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4391_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_51_2 ), .O(n5774));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4391_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13415_bdd_4_lut (.I0(n13415), .I1(\REG.mem_53_13 ), .I2(\REG.mem_52_13 ), 
            .I3(rd_addr_r_c[1]), .O(n13418));
    defparam n13415_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10597 (.I0(rd_addr_r_c[1]), .I1(n11246), 
            .I2(n11247), .I3(rd_addr_r_c[2]), .O(n12305));
    defparam rd_addr_r_1__bdd_4_lut_10597.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10568 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_13 ), 
            .I2(\REG.mem_3_13 ), .I3(rd_addr_r_c[1]), .O(n12425));
    defparam rd_addr_r_0__bdd_4_lut_10568.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11385 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_6 ), 
            .I2(\REG.mem_59_6 ), .I3(rd_addr_r_c[1]), .O(n13409));
    defparam rd_addr_r_0__bdd_4_lut_11385.LUT_INIT = 16'he4aa;
    SB_DFF i245_246 (.Q(\REG.mem_2_5 ), .C(FIFO_CLK_c), .D(n4950));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13409_bdd_4_lut (.I0(n13409), .I1(\REG.mem_57_6 ), .I2(\REG.mem_56_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11593));
    defparam n13409_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4390_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_51_1 ), .O(n5773));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4390_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10846 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_11 ), 
            .I2(\REG.mem_63_11 ), .I3(rd_addr_r_c[1]), .O(n12761));
    defparam rd_addr_r_0__bdd_4_lut_10846.LUT_INIT = 16'he4aa;
    SB_LUT4 i4389_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_51_0 ), .O(n5772));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4389_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12761_bdd_4_lut (.I0(n12761), .I1(\REG.mem_61_11 ), .I2(\REG.mem_60_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11737));
    defparam n12761_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4093_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_34_1 ), .O(n5476));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4093_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9194_3_lut (.I0(n12698), .I1(n13802), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [2]));
    defparam i9194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9437_3_lut (.I0(n12884), .I1(n13160), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [4]));
    defparam i9437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9689_3_lut (.I0(n13028), .I1(n13586), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [5]));
    defparam i9689_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR full_ext_r_117 (.Q(full_o), .C(FIFO_CLK_c), .D(full_nxt_c_N_626), 
            .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 i9553_3_lut (.I0(n12992), .I1(n12824), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11391));
    defparam i9553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9554_3_lut (.I0(n12962), .I1(n11391), .I2(rd_addr_r_c[3]), 
            .I3(GND_net), .O(n11392));
    defparam i9554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11390 (.I0(rd_addr_r_c[1]), .I1(n11531), 
            .I2(n11532), .I3(rd_addr_r_c[2]), .O(n13403));
    defparam rd_addr_r_1__bdd_4_lut_11390.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10841 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_0 ), 
            .I2(\REG.mem_35_0 ), .I3(rd_addr_r_c[1]), .O(n12755));
    defparam rd_addr_r_0__bdd_4_lut_10841.LUT_INIT = 16'he4aa;
    SB_DFFE \REG.out_raw__i1  (.Q(\REG.out_raw[0] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [0]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_LUT4 i9779_3_lut (.I0(n13088), .I1(n13334), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [7]));
    defparam i9779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13403_bdd_4_lut (.I0(n13403), .I1(n11511), .I2(n11510), .I3(rd_addr_r_c[2]), 
            .O(n11595));
    defparam n13403_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9260_3_lut (.I0(n12788), .I1(n13286), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [8]));
    defparam i9260_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i242_243 (.Q(\REG.mem_2_4 ), .C(FIFO_CLK_c), .D(n4949));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9764_3_lut (.I0(n13082), .I1(n13376), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [10]));
    defparam i9764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12755_bdd_4_lut (.I0(n12755), .I1(\REG.mem_33_0 ), .I2(\REG.mem_32_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11320));
    defparam n12755_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9682_3_lut (.I0(\REG.mem_54_10 ), .I1(\REG.mem_55_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11520));
    defparam i9682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i76_2_lut_3_lut_4_lut (.I0(n20_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n62));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i76_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i9681_3_lut (.I0(\REG.mem_52_10 ), .I1(\REG.mem_53_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11519));
    defparam i9681_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i239_240 (.Q(\REG.mem_2_3 ), .C(FIFO_CLK_c), .D(n4948));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i75_2_lut_3_lut_4_lut (.I0(n20_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n30));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i75_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11380 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_3 ), 
            .I2(\REG.mem_31_3 ), .I3(rd_addr_r_c[1]), .O(n13397));
    defparam rd_addr_r_0__bdd_4_lut_11380.LUT_INIT = 16'he4aa;
    SB_LUT4 i10097_3_lut (.I0(n13484), .I1(n13748), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [12]));
    defparam i10097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9278_3_lut (.I0(n12800), .I1(n13238), .I2(rd_addr_r_c[3]), 
            .I3(GND_net), .O(n11116));
    defparam i9278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9346_3_lut (.I0(n11116), .I1(n12638), .I2(rd_addr_r_c[4]), 
            .I3(GND_net), .O(n11184));
    defparam i9346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13397_bdd_4_lut (.I0(n13397), .I1(\REG.mem_29_3 ), .I2(\REG.mem_28_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11077));
    defparam n13397_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9347_3_lut (.I0(n12842), .I1(n11184), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [14]));
    defparam i9347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9224_3_lut (.I0(n12734), .I1(n13532), .I2(rd_addr_r_c[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [15]));
    defparam i9224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9636_3_lut (.I0(\REG.mem_48_7 ), .I1(\REG.mem_49_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11474));
    defparam i9636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9637_3_lut (.I0(\REG.mem_50_7 ), .I1(\REG.mem_51_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11475));
    defparam i9637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9667_3_lut (.I0(\REG.mem_54_7 ), .I1(\REG.mem_55_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11505));
    defparam i9667_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i236_237 (.Q(\REG.mem_2_2 ), .C(FIFO_CLK_c), .D(n4947));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9666_3_lut (.I0(\REG.mem_52_7 ), .I1(\REG.mem_53_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11504));
    defparam i9666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10866 (.I0(rd_addr_r_c[2]), .I1(n11068), 
            .I2(n11077), .I3(rd_addr_r_c[3]), .O(n12749));
    defparam rd_addr_r_2__bdd_4_lut_10866.LUT_INIT = 16'he4aa;
    SB_LUT4 i4091_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_34_0 ), .O(n5474));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4091_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12425_bdd_4_lut (.I0(n12425), .I1(\REG.mem_1_13 ), .I2(\REG.mem_0_13 ), 
            .I3(rd_addr_r_c[1]), .O(n11815));
    defparam n12425_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12749_bdd_4_lut (.I0(n12749), .I1(n11065), .I2(n11059), .I3(rd_addr_r_c[3]), 
            .O(n11137));
    defparam n12749_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11375 (.I0(rd_addr_r_c[1]), .I1(n11555), 
            .I2(n11556), .I3(rd_addr_r_c[2]), .O(n13391));
    defparam rd_addr_r_1__bdd_4_lut_11375.LUT_INIT = 16'he4aa;
    SB_LUT4 i9678_3_lut (.I0(\REG.mem_48_10 ), .I1(\REG.mem_49_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11516));
    defparam i9678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9679_3_lut (.I0(\REG.mem_50_10 ), .I1(\REG.mem_51_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11517));
    defparam i9679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10871 (.I0(rd_addr_r_c[1]), .I1(n11870), 
            .I2(n11871), .I3(rd_addr_r_c[2]), .O(n12743));
    defparam rd_addr_r_1__bdd_4_lut_10871.LUT_INIT = 16'he4aa;
    SB_LUT4 n13391_bdd_4_lut (.I0(n13391), .I1(n11541), .I2(n11540), .I3(rd_addr_r_c[2]), 
            .O(n13394));
    defparam n13391_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i6_2_lut_4_lut (.I0(wr_grey_sync_r[6]), 
            .I1(wr_addr_p1_w[6]), .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[5] ), 
            .O(wr_grey_w[5]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i6_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 n12743_bdd_4_lut (.I0(n12743), .I1(n11868), .I2(n11867), .I3(rd_addr_r_c[2]), 
            .O(n12746));
    defparam n12743_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9604_3_lut (.I0(\REG.mem_22_8 ), .I1(\REG.mem_23_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11442));
    defparam i9604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10563 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_9 ), 
            .I2(\REG.mem_59_9 ), .I3(rd_addr_r_c[1]), .O(n12419));
    defparam rd_addr_r_0__bdd_4_lut_10563.LUT_INIT = 16'he4aa;
    SB_LUT4 i9603_3_lut (.I0(\REG.mem_20_8 ), .I1(\REG.mem_21_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11441));
    defparam i9603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11370 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_5 ), 
            .I2(\REG.mem_27_5 ), .I3(rd_addr_r_c[1]), .O(n13385));
    defparam rd_addr_r_0__bdd_4_lut_11370.LUT_INIT = 16'he4aa;
    SB_LUT4 i4289_2_lut_4_lut (.I0(wr_grey_sync_r[6]), .I1(wr_addr_p1_w[6]), 
            .I2(wr_sig_mv_w), .I3(reset_per_frame), .O(n5672));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i4289_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 n13385_bdd_4_lut (.I0(n13385), .I1(\REG.mem_25_5 ), .I2(\REG.mem_24_5 ), 
            .I3(rd_addr_r_c[1]), .O(n13388));
    defparam n13385_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR rd_grey_sync_r__i0 (.Q(\rd_grey_sync_r[0] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[0]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10836 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_15 ), 
            .I2(\REG.mem_27_15 ), .I3(rd_addr_r_c[1]), .O(n12737));
    defparam rd_addr_r_0__bdd_4_lut_10836.LUT_INIT = 16'he4aa;
    SB_LUT4 n12737_bdd_4_lut (.I0(n12737), .I1(\REG.mem_25_15 ), .I2(\REG.mem_24_15 ), 
            .I3(rd_addr_r_c[1]), .O(n12740));
    defparam n12737_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9730_3_lut (.I0(n12326), .I1(n13850), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11568));
    defparam i9730_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i233_234 (.Q(\REG.mem_2_1 ), .C(FIFO_CLK_c), .D(n4946));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9729_3_lut (.I0(n12542), .I1(n12362), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11567));
    defparam i9729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11360 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_12 ), 
            .I2(\REG.mem_15_12 ), .I3(rd_addr_r_c[1]), .O(n13379));
    defparam rd_addr_r_0__bdd_4_lut_11360.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10861 (.I0(rd_addr_r_c[3]), .I1(n12650), 
            .I2(n11016), .I3(rd_addr_r_c[4]), .O(n12731));
    defparam rd_addr_r_3__bdd_4_lut_10861.LUT_INIT = 16'he4aa;
    SB_DFFSS empty_ext_r_124 (.Q(DEBUG_3_c), .C(SLM_CLK_c), .D(empty_nxt_c_N_629), 
            .S(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_LUT4 n13379_bdd_4_lut (.I0(n13379), .I1(\REG.mem_13_12 ), .I2(\REG.mem_12_12 ), 
            .I3(rd_addr_r_c[1]), .O(n13382));
    defparam n13379_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i230_231 (.Q(\REG.mem_2_0 ), .C(FIFO_CLK_c), .D(n4945));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFSR wr_grey_sync_r__i0 (.Q(wr_grey_sync_r[0]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[0]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFF i38_39 (.Q(\REG.mem_0_0 ), .C(FIFO_CLK_c), .D(n4944));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11440 (.I0(rd_addr_r_c[3]), .I1(n13070), 
            .I2(n11586), .I3(rd_addr_r_c[4]), .O(n13373));
    defparam rd_addr_r_3__bdd_4_lut_11440.LUT_INIT = 16'he4aa;
    SB_DFF i41_42 (.Q(\REG.mem_0_1 ), .C(FIFO_CLK_c), .D(n4943));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFS \aempty_flag_impl.ae_flag_ext_r_130  (.Q(dc32_fifo_almost_empty), 
            .C(SLM_CLK_c), .D(\aempty_flag_impl.ae_flag_nxt_w ), .S(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(669[37] 672[40])
    SB_LUT4 i9715_3_lut (.I0(n13154), .I1(n12656), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11553));
    defparam i9715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12731_bdd_4_lut (.I0(n12731), .I1(n11952), .I2(n11951), .I3(rd_addr_r_c[4]), 
            .O(n12734));
    defparam n12731_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13373_bdd_4_lut (.I0(n13373), .I1(n11562), .I2(n13052), .I3(rd_addr_r_c[4]), 
            .O(n13376));
    defparam n13373_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11355 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_1 ), 
            .I2(\REG.mem_7_1 ), .I3(rd_addr_r_c[1]), .O(n13367));
    defparam rd_addr_r_0__bdd_4_lut_11355.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10831 (.I0(rd_addr_r_c[2]), .I1(n11623), 
            .I2(n11632), .I3(rd_addr_r_c[3]), .O(n12725));
    defparam rd_addr_r_2__bdd_4_lut_10831.LUT_INIT = 16'he4aa;
    SB_LUT4 n13367_bdd_4_lut (.I0(n13367), .I1(\REG.mem_5_1 ), .I2(\REG.mem_4_1 ), 
            .I3(rd_addr_r_c[1]), .O(n11230));
    defparam n13367_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12419_bdd_4_lut (.I0(n12419), .I1(\REG.mem_57_9 ), .I2(\REG.mem_56_9 ), 
            .I3(rd_addr_r_c[1]), .O(n12422));
    defparam n12419_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12725_bdd_4_lut (.I0(n12725), .I1(n11611), .I2(n11608), .I3(rd_addr_r_c[3]), 
            .O(n11743));
    defparam n12725_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9181_3_lut (.I0(n13778), .I1(n13754), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11019));
    defparam i9181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10826 (.I0(rd_addr_r_c[1]), .I1(n11894), 
            .I2(n11895), .I3(rd_addr_r_c[2]), .O(n12719));
    defparam rd_addr_r_1__bdd_4_lut_10826.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11345 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_3 ), 
            .I2(\REG.mem_35_3 ), .I3(rd_addr_r_c[1]), .O(n13361));
    defparam rd_addr_r_0__bdd_4_lut_11345.LUT_INIT = 16'he4aa;
    SB_LUT4 n13361_bdd_4_lut (.I0(n13361), .I1(\REG.mem_33_3 ), .I2(\REG.mem_32_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11080));
    defparam n13361_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12719_bdd_4_lut (.I0(n12719), .I1(n11883), .I2(n11882), .I3(rd_addr_r_c[2]), 
            .O(n12722));
    defparam n12719_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11340 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_1 ), 
            .I2(\REG.mem_47_1 ), .I3(rd_addr_r_c[1]), .O(n13355));
    defparam rd_addr_r_0__bdd_4_lut_11340.LUT_INIT = 16'he4aa;
    SB_LUT4 n13355_bdd_4_lut (.I0(n13355), .I1(\REG.mem_45_1 ), .I2(\REG.mem_44_1 ), 
            .I3(rd_addr_r_c[1]), .O(n13358));
    defparam n13355_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10047_3_lut (.I0(\REG.mem_24_2 ), .I1(\REG.mem_25_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11885));
    defparam i10047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10806 (.I0(rd_addr_r_c[1]), .I1(n11864), 
            .I2(n11865), .I3(rd_addr_r_c[2]), .O(n12713));
    defparam rd_addr_r_1__bdd_4_lut_10806.LUT_INIT = 16'he4aa;
    SB_LUT4 i3825_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_17_15 ), .O(n5208));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3825_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3824_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_17_14 ), .O(n5207));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3824_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10048_3_lut (.I0(\REG.mem_26_2 ), .I1(\REG.mem_27_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11886));
    defparam i10048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3823_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_17_13 ), .O(n5206));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3823_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11335 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_11 ), 
            .I2(\REG.mem_3_11 ), .I3(rd_addr_r_c[1]), .O(n13349));
    defparam rd_addr_r_0__bdd_4_lut_11335.LUT_INIT = 16'he4aa;
    SB_DFF i44_45 (.Q(\REG.mem_0_2 ), .C(FIFO_CLK_c), .D(n4941));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13349_bdd_4_lut (.I0(n13349), .I1(\REG.mem_1_11 ), .I2(\REG.mem_0_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11608));
    defparam n13349_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12713_bdd_4_lut (.I0(n12713), .I1(n11856), .I2(n11855), .I3(rd_addr_r_c[2]), 
            .O(n12716));
    defparam n12713_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10060_3_lut (.I0(\REG.mem_30_2 ), .I1(\REG.mem_31_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11898));
    defparam i10060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10059_3_lut (.I0(\REG.mem_28_2 ), .I1(\REG.mem_29_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11897));
    defparam i10059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10821 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_12 ), 
            .I2(\REG.mem_51_12 ), .I3(rd_addr_r_c[1]), .O(n12707));
    defparam rd_addr_r_0__bdd_4_lut_10821.LUT_INIT = 16'he4aa;
    SB_LUT4 i3822_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_17_12 ), .O(n5205));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3822_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11330 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_11 ), 
            .I2(\REG.mem_7_11 ), .I3(rd_addr_r_c[1]), .O(n13343));
    defparam rd_addr_r_0__bdd_4_lut_11330.LUT_INIT = 16'he4aa;
    SB_LUT4 n13343_bdd_4_lut (.I0(n13343), .I1(\REG.mem_5_11 ), .I2(\REG.mem_4_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11611));
    defparam n13343_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3821_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_17_11 ), .O(n5204));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3821_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12305_bdd_4_lut (.I0(n12305), .I1(n11232), .I2(n11231), .I3(rd_addr_r_c[2]), 
            .O(n12308));
    defparam n12305_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12707_bdd_4_lut (.I0(n12707), .I1(\REG.mem_49_12 ), .I2(\REG.mem_48_12 ), 
            .I3(rd_addr_r_c[1]), .O(n12710));
    defparam n12707_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10474 (.I0(rd_addr_r_c[2]), .I1(n11965), 
            .I2(n11971), .I3(rd_addr_r_c[3]), .O(n12311));
    defparam rd_addr_r_2__bdd_4_lut_10474.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10479 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_4 ), 
            .I2(\REG.mem_3_4 ), .I3(rd_addr_r_c[1]), .O(n12299));
    defparam rd_addr_r_0__bdd_4_lut_10479.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10796 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_8 ), 
            .I2(\REG.mem_15_8 ), .I3(rd_addr_r_c[1]), .O(n12701));
    defparam rd_addr_r_0__bdd_4_lut_10796.LUT_INIT = 16'he4aa;
    SB_LUT4 i10020_3_lut (.I0(\REG.mem_8_14 ), .I1(\REG.mem_9_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11858));
    defparam i10020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3820_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_17_10 ), .O(n5203));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3820_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10021_3_lut (.I0(\REG.mem_10_14 ), .I1(\REG.mem_11_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11859));
    defparam i10021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11325 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_6 ), 
            .I2(\REG.mem_63_6 ), .I3(rd_addr_r_c[1]), .O(n13337));
    defparam rd_addr_r_0__bdd_4_lut_11325.LUT_INIT = 16'he4aa;
    SB_DFF i47_48 (.Q(\REG.mem_0_3 ), .C(FIFO_CLK_c), .D(n4940));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12701_bdd_4_lut (.I0(n12701), .I1(\REG.mem_13_8 ), .I2(\REG.mem_12_8 ), 
            .I3(rd_addr_r_c[1]), .O(n12704));
    defparam n12701_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10024_3_lut (.I0(\REG.mem_14_14 ), .I1(\REG.mem_15_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11862));
    defparam i10024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10816 (.I0(rd_addr_r_c[3]), .I1(n11012), 
            .I2(n12470), .I3(rd_addr_r_c[4]), .O(n12695));
    defparam rd_addr_r_3__bdd_4_lut_10816.LUT_INIT = 16'he4aa;
    SB_LUT4 i3819_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_17_9 ), .O(n5202));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3819_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3818_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_17_8 ), .O(n5201));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3818_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10558 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_1 ), 
            .I2(\REG.mem_3_1 ), .I3(rd_addr_r_c[1]), .O(n12413));
    defparam rd_addr_r_0__bdd_4_lut_10558.LUT_INIT = 16'he4aa;
    SB_LUT4 i3817_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_17_7 ), .O(n5200));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3817_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12695_bdd_4_lut (.I0(n12695), .I1(n11010), .I2(n11009), .I3(rd_addr_r_c[4]), 
            .O(n12698));
    defparam n12695_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10023_3_lut (.I0(\REG.mem_12_14 ), .I1(\REG.mem_13_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11861));
    defparam i10023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10801 (.I0(rd_addr_r_c[1]), .I1(n11852), 
            .I2(n11853), .I3(rd_addr_r_c[2]), .O(n12689));
    defparam rd_addr_r_1__bdd_4_lut_10801.LUT_INIT = 16'he4aa;
    SB_LUT4 n13337_bdd_4_lut (.I0(n13337), .I1(\REG.mem_61_6 ), .I2(\REG.mem_60_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11614));
    defparam n13337_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3816_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_17_6 ), .O(n5199));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3816_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12689_bdd_4_lut (.I0(n12689), .I1(n11850), .I2(n11849), .I3(rd_addr_r_c[2]), 
            .O(n12692));
    defparam n12689_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3815_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_17_5 ), .O(n5198));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3815_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3814_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_17_4 ), .O(n5197));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3814_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11350 (.I0(rd_addr_r_c[3]), .I1(n13076), 
            .I2(n11595), .I3(rd_addr_r_c[4]), .O(n13331));
    defparam rd_addr_r_3__bdd_4_lut_11350.LUT_INIT = 16'he4aa;
    SB_LUT4 n13331_bdd_4_lut (.I0(n13331), .I1(n11583), .I2(n13064), .I3(rd_addr_r_c[4]), 
            .O(n13334));
    defparam n13331_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3813_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_17_3 ), .O(n5196));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3813_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10791 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_8 ), 
            .I2(\REG.mem_43_8 ), .I3(rd_addr_r_c[1]), .O(n12683));
    defparam rd_addr_r_0__bdd_4_lut_10791.LUT_INIT = 16'he4aa;
    SB_LUT4 i3812_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_17_2 ), .O(n5195));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3812_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3811_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_17_1 ), .O(n5194));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3811_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11365 (.I0(rd_addr_r_c[1]), .I1(n11171), 
            .I2(n11172), .I3(rd_addr_r_c[2]), .O(n13325));
    defparam rd_addr_r_1__bdd_4_lut_11365.LUT_INIT = 16'he4aa;
    SB_LUT4 n13325_bdd_4_lut (.I0(n13325), .I1(n11169), .I2(n11168), .I3(rd_addr_r_c[2]), 
            .O(n11250));
    defparam n13325_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12683_bdd_4_lut (.I0(n12683), .I1(\REG.mem_41_8 ), .I2(\REG.mem_40_8 ), 
            .I3(rd_addr_r_c[1]), .O(n12686));
    defparam n12683_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3810_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_17_0 ), .O(n5193));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3810_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_addr_r_6__I_0_135_i6_3_lut (.I0(wr_addr_r[5]), .I1(wr_addr_p1_w[5]), 
            .I2(wr_sig_mv_w), .I3(GND_net), .O(\wr_addr_nxt_c[5] ));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_6__I_0_135_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10782 (.I0(rd_addr_r_c[1]), .I1(n11948), 
            .I2(n11949), .I3(rd_addr_r_c[2]), .O(n12677));
    defparam rd_addr_r_1__bdd_4_lut_10782.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11320 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_12 ), 
            .I2(\REG.mem_19_12 ), .I3(rd_addr_r_c[1]), .O(n13319));
    defparam rd_addr_r_0__bdd_4_lut_11320.LUT_INIT = 16'he4aa;
    SB_LUT4 n12413_bdd_4_lut (.I0(n12413), .I1(\REG.mem_1_1 ), .I2(\REG.mem_0_1 ), 
            .I3(rd_addr_r_c[1]), .O(n12416));
    defparam n12413_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3857_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_19_15 ), .O(n5240));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3857_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13319_bdd_4_lut (.I0(n13319), .I1(\REG.mem_17_12 ), .I2(\REG.mem_16_12 ), 
            .I3(rd_addr_r_c[1]), .O(n13322));
    defparam n13319_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3856_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_19_14 ), .O(n5239));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3856_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3855_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_19_13 ), .O(n5238));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3855_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12677_bdd_4_lut (.I0(n12677), .I1(n11943), .I2(n11942), .I3(rd_addr_r_c[2]), 
            .O(n12680));
    defparam n12677_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3854_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_19_12 ), .O(n5237));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3854_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3853_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_19_11 ), .O(n5236));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3853_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3852_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_19_10 ), .O(n5235));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3852_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3851_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_19_9 ), .O(n5234));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3851_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3850_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_19_8 ), .O(n5233));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3850_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10772 (.I0(rd_addr_r_c[1]), .I1(n11909), 
            .I2(n11910), .I3(rd_addr_r_c[2]), .O(n12671));
    defparam rd_addr_r_1__bdd_4_lut_10772.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11310 (.I0(rd_addr_r_c[1]), .I1(n11198), 
            .I2(n11199), .I3(rd_addr_r_c[2]), .O(n13313));
    defparam rd_addr_r_1__bdd_4_lut_11310.LUT_INIT = 16'he4aa;
    SB_LUT4 i3849_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_19_7 ), .O(n5232));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3849_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12671_bdd_4_lut (.I0(n12671), .I1(n11907), .I2(n11906), .I3(rd_addr_r_c[2]), 
            .O(n12674));
    defparam n12671_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3848_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_19_6 ), .O(n5231));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3848_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10777 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_15 ), 
            .I2(\REG.mem_31_15 ), .I3(rd_addr_r_c[1]), .O(n12665));
    defparam rd_addr_r_0__bdd_4_lut_10777.LUT_INIT = 16'he4aa;
    SB_LUT4 n13313_bdd_4_lut (.I0(n13313), .I1(n11193), .I2(n11192), .I3(rd_addr_r_c[2]), 
            .O(n11256));
    defparam n13313_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3847_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_19_5 ), .O(n5230));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3847_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3846_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_19_4 ), .O(n5229));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3846_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3845_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_19_3 ), .O(n5228));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3845_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12665_bdd_4_lut (.I0(n12665), .I1(\REG.mem_29_15 ), .I2(\REG.mem_28_15 ), 
            .I3(rd_addr_r_c[1]), .O(n12668));
    defparam n12665_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11305 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_3 ), 
            .I2(\REG.mem_39_3 ), .I3(rd_addr_r_c[1]), .O(n13307));
    defparam rd_addr_r_0__bdd_4_lut_11305.LUT_INIT = 16'he4aa;
    SB_LUT4 n13307_bdd_4_lut (.I0(n13307), .I1(\REG.mem_37_3 ), .I2(\REG.mem_36_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11086));
    defparam n13307_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10811 (.I0(rd_addr_r_c[2]), .I1(n11656), 
            .I2(n11668), .I3(rd_addr_r_c[3]), .O(n12659));
    defparam rd_addr_r_2__bdd_4_lut_10811.LUT_INIT = 16'he4aa;
    SB_LUT4 n12659_bdd_4_lut (.I0(n12659), .I1(n11653), .I2(n11644), .I3(rd_addr_r_c[3]), 
            .O(n11755));
    defparam n12659_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3844_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_19_2 ), .O(n5227));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3844_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11295 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_3 ), 
            .I2(\REG.mem_43_3 ), .I3(rd_addr_r_c[1]), .O(n13301));
    defparam rd_addr_r_0__bdd_4_lut_11295.LUT_INIT = 16'he4aa;
    SB_LUT4 i3843_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_19_1 ), .O(n5226));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3843_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10762 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_7 ), 
            .I2(\REG.mem_15_7 ), .I3(rd_addr_r_c[1]), .O(n12653));
    defparam rd_addr_r_0__bdd_4_lut_10762.LUT_INIT = 16'he4aa;
    SB_LUT4 n12653_bdd_4_lut (.I0(n12653), .I1(\REG.mem_13_7 ), .I2(\REG.mem_12_7 ), 
            .I3(rd_addr_r_c[1]), .O(n12656));
    defparam n12653_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13301_bdd_4_lut (.I0(n13301), .I1(\REG.mem_41_3 ), .I2(\REG.mem_40_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11089));
    defparam n13301_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10767 (.I0(rd_addr_r_c[1]), .I1(n11714), 
            .I2(n11715), .I3(rd_addr_r_c[2]), .O(n12647));
    defparam rd_addr_r_1__bdd_4_lut_10767.LUT_INIT = 16'he4aa;
    SB_LUT4 i3842_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_19_0 ), .O(n5225));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3842_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12647_bdd_4_lut (.I0(n12647), .I1(n11694), .I2(n11693), .I3(rd_addr_r_c[2]), 
            .O(n12650));
    defparam n12647_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11290 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_0 ), 
            .I2(\REG.mem_59_0 ), .I3(rd_addr_r_c[1]), .O(n13295));
    defparam rd_addr_r_0__bdd_4_lut_11290.LUT_INIT = 16'he4aa;
    SB_LUT4 n13295_bdd_4_lut (.I0(n13295), .I1(\REG.mem_57_0 ), .I2(\REG.mem_56_0 ), 
            .I3(rd_addr_r_c[1]), .O(n13298));
    defparam n13295_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10747 (.I0(rd_addr_r_c[1]), .I1(n11681), 
            .I2(n11682), .I3(rd_addr_r_c[2]), .O(n12641));
    defparam rd_addr_r_1__bdd_4_lut_10747.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11285 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_11 ), 
            .I2(\REG.mem_11_11 ), .I3(rd_addr_r_c[1]), .O(n13289));
    defparam rd_addr_r_0__bdd_4_lut_11285.LUT_INIT = 16'he4aa;
    SB_LUT4 n12641_bdd_4_lut (.I0(n12641), .I1(n11637), .I2(n11636), .I3(rd_addr_r_c[2]), 
            .O(n12644));
    defparam n12641_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13289_bdd_4_lut (.I0(n13289), .I1(\REG.mem_9_11 ), .I2(\REG.mem_8_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11623));
    defparam n13289_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10553 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_12 ), 
            .I2(\REG.mem_63_12 ), .I3(rd_addr_r_c[1]), .O(n12407));
    defparam rd_addr_r_0__bdd_4_lut_10553.LUT_INIT = 16'he4aa;
    SB_LUT4 i3873_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_20_15 ), .O(n5256));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3873_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3872_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_20_14 ), .O(n5255));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3872_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3871_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_20_13 ), .O(n5254));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3871_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3870_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_20_12 ), .O(n5253));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3870_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3869_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_20_11 ), .O(n5252));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3869_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3868_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_20_10 ), .O(n5251));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3868_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10757 (.I0(rd_addr_r_c[2]), .I1(n10993), 
            .I2(n10996), .I3(rd_addr_r_c[3]), .O(n12635));
    defparam rd_addr_r_2__bdd_4_lut_10757.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11315 (.I0(rd_addr_r_c[3]), .I1(n12716), 
            .I2(n11049), .I3(rd_addr_r_c[4]), .O(n13283));
    defparam rd_addr_r_3__bdd_4_lut_11315.LUT_INIT = 16'he4aa;
    SB_LUT4 n12635_bdd_4_lut (.I0(n12635), .I1(n12016), .I2(n12010), .I3(rd_addr_r_c[3]), 
            .O(n12638));
    defparam n12635_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3867_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_20_9 ), .O(n5250));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3867_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10752 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_12 ), 
            .I2(\REG.mem_55_12 ), .I3(rd_addr_r_c[1]), .O(n12629));
    defparam rd_addr_r_0__bdd_4_lut_10752.LUT_INIT = 16'he4aa;
    SB_LUT4 n13283_bdd_4_lut (.I0(n13283), .I1(n11004), .I2(n12644), .I3(rd_addr_r_c[4]), 
            .O(n13286));
    defparam n13283_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12629_bdd_4_lut (.I0(n12629), .I1(\REG.mem_53_12 ), .I2(\REG.mem_52_12 ), 
            .I3(rd_addr_r_c[1]), .O(n12632));
    defparam n12629_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11300 (.I0(rd_addr_r_c[1]), .I1(n11219), 
            .I2(n11220), .I3(rd_addr_r_c[2]), .O(n13277));
    defparam rd_addr_r_1__bdd_4_lut_11300.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10732 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_15 ), 
            .I2(\REG.mem_35_15 ), .I3(rd_addr_r_c[1]), .O(n12623));
    defparam rd_addr_r_0__bdd_4_lut_10732.LUT_INIT = 16'he4aa;
    SB_LUT4 n12623_bdd_4_lut (.I0(n12623), .I1(\REG.mem_33_15 ), .I2(\REG.mem_32_15 ), 
            .I3(rd_addr_r_c[1]), .O(n12626));
    defparam n12623_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13277_bdd_4_lut (.I0(n13277), .I1(n11217), .I2(n11216), .I3(rd_addr_r_c[2]), 
            .O(n11259));
    defparam n13277_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11280 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_15 ), 
            .I2(\REG.mem_3_15 ), .I3(rd_addr_r_c[1]), .O(n13271));
    defparam rd_addr_r_0__bdd_4_lut_11280.LUT_INIT = 16'he4aa;
    SB_LUT4 i3866_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_20_8 ), .O(n5249));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3866_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3865_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_20_7 ), .O(n5248));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3865_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_addr_r_6__I_0_135_i4_3_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_w[3]), 
            .I2(wr_sig_mv_w), .I3(GND_net), .O(\wr_addr_nxt_c[3] ));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_6__I_0_135_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13271_bdd_4_lut (.I0(n13271), .I1(\REG.mem_1_15 ), .I2(\REG.mem_0_15 ), 
            .I3(rd_addr_r_c[1]), .O(n13274));
    defparam n13271_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i50_51 (.Q(\REG.mem_0_4 ), .C(FIFO_CLK_c), .D(n4935));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10727 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_9 ), 
            .I2(\REG.mem_51_9 ), .I3(rd_addr_r_c[1]), .O(n12617));
    defparam rd_addr_r_0__bdd_4_lut_10727.LUT_INIT = 16'he4aa;
    SB_DFF i53_54 (.Q(\REG.mem_0_5 ), .C(FIFO_CLK_c), .D(n4934));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12617_bdd_4_lut (.I0(n12617), .I1(\REG.mem_49_9 ), .I2(\REG.mem_48_9 ), 
            .I3(rd_addr_r_c[1]), .O(n12620));
    defparam n12617_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3864_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_20_6 ), .O(n5247));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3864_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3863_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_20_5 ), .O(n5246));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3863_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12299_bdd_4_lut (.I0(n12299), .I1(\REG.mem_1_4 ), .I2(\REG.mem_0_4 ), 
            .I3(rd_addr_r_c[1]), .O(n12302));
    defparam n12299_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10460 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_8 ), 
            .I2(\REG.mem_47_8 ), .I3(rd_addr_r_c[1]), .O(n12293));
    defparam rd_addr_r_0__bdd_4_lut_10460.LUT_INIT = 16'he4aa;
    SB_LUT4 i3862_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_20_4 ), .O(n5245));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3862_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3861_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_20_3 ), .O(n5244));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3861_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11265 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_3 ), 
            .I2(\REG.mem_47_3 ), .I3(rd_addr_r_c[1]), .O(n13265));
    defparam rd_addr_r_0__bdd_4_lut_11265.LUT_INIT = 16'he4aa;
    SB_LUT4 n12293_bdd_4_lut (.I0(n12293), .I1(\REG.mem_45_8 ), .I2(\REG.mem_44_8 ), 
            .I3(rd_addr_r_c[1]), .O(n12296));
    defparam n12293_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12335_bdd_4_lut (.I0(n12335), .I1(\REG.mem_17_2 ), .I2(\REG.mem_16_2 ), 
            .I3(rd_addr_r_c[1]), .O(n12338));
    defparam n12335_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10489 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_9 ), 
            .I2(\REG.mem_11_9 ), .I3(rd_addr_r_c[1]), .O(n12329));
    defparam rd_addr_r_0__bdd_4_lut_10489.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10737 (.I0(rd_addr_r_c[2]), .I1(n11692), 
            .I2(n11701), .I3(rd_addr_r_c[3]), .O(n12611));
    defparam rd_addr_r_2__bdd_4_lut_10737.LUT_INIT = 16'he4aa;
    SB_LUT4 n13265_bdd_4_lut (.I0(n13265), .I1(\REG.mem_45_3 ), .I2(\REG.mem_44_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11104));
    defparam n13265_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3860_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_20_2 ), .O(n5243));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3860_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3859_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_20_1 ), .O(n5242));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3859_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12323_bdd_4_lut (.I0(n12323), .I1(\REG.mem_25_7 ), .I2(\REG.mem_24_7 ), 
            .I3(rd_addr_r_c[1]), .O(n12326));
    defparam n12323_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11260 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_12 ), 
            .I2(\REG.mem_23_12 ), .I3(rd_addr_r_c[1]), .O(n13259));
    defparam rd_addr_r_0__bdd_4_lut_11260.LUT_INIT = 16'he4aa;
    SB_LUT4 i3858_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_20_0 ), .O(n5241));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3858_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12611_bdd_4_lut (.I0(n12611), .I1(n11677), .I2(n11674), .I3(rd_addr_r_c[3]), 
            .O(n11764));
    defparam n12611_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10587 (.I0(rd_addr_r_c[2]), .I1(n11158), 
            .I2(n11176), .I3(rd_addr_r_c[3]), .O(n12317));
    defparam rd_addr_r_2__bdd_4_lut_10587.LUT_INIT = 16'he4aa;
    SB_LUT4 i3890_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_21_15 ), .O(n5273));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3890_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13259_bdd_4_lut (.I0(n13259), .I1(\REG.mem_21_12 ), .I2(\REG.mem_20_12 ), 
            .I3(rd_addr_r_c[1]), .O(n13262));
    defparam n13259_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12407_bdd_4_lut (.I0(n12407), .I1(\REG.mem_61_12 ), .I2(\REG.mem_60_12 ), 
            .I3(rd_addr_r_c[1]), .O(n12410));
    defparam n12407_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12311_bdd_4_lut (.I0(n12311), .I1(n11959), .I2(n11815), .I3(rd_addr_r_c[3]), 
            .O(n12314));
    defparam n12311_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3889_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_21_14 ), .O(n5272));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3889_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3888_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_21_13 ), .O(n5271));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3888_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10494 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_2 ), 
            .I2(\REG.mem_19_2 ), .I3(rd_addr_r_c[1]), .O(n12335));
    defparam rd_addr_r_0__bdd_4_lut_10494.LUT_INIT = 16'he4aa;
    SB_LUT4 i3887_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_21_12 ), .O(n5270));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3887_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3886_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_21_11 ), .O(n5269));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3886_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i5_1_lut (.I0(rd_addr_r_c[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3885_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_21_10 ), .O(n5268));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3885_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3884_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_21_9 ), .O(n5267));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3884_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10722 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_0 ), 
            .I2(\REG.mem_39_0 ), .I3(rd_addr_r_c[1]), .O(n12605));
    defparam rd_addr_r_0__bdd_4_lut_10722.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10469 (.I0(rd_addr_r_c[2]), .I1(n11455), 
            .I2(n11488), .I3(rd_addr_r_c[3]), .O(n12287));
    defparam rd_addr_r_2__bdd_4_lut_10469.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11255 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_13 ), 
            .I2(\REG.mem_31_13 ), .I3(rd_addr_r_c[1]), .O(n13253));
    defparam rd_addr_r_0__bdd_4_lut_11255.LUT_INIT = 16'he4aa;
    SB_LUT4 n12605_bdd_4_lut (.I0(n12605), .I1(\REG.mem_37_0 ), .I2(\REG.mem_36_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11332));
    defparam n12605_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13253_bdd_4_lut (.I0(n13253), .I1(\REG.mem_29_13 ), .I2(\REG.mem_28_13 ), 
            .I3(rd_addr_r_c[1]), .O(n13256));
    defparam n13253_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3883_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_21_8 ), .O(n5266));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3883_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10717 (.I0(rd_addr_r_c[2]), .I1(n11722), 
            .I2(n11737), .I3(rd_addr_r_c[3]), .O(n12599));
    defparam rd_addr_r_2__bdd_4_lut_10717.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11250 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_6 ), 
            .I2(\REG.mem_19_6 ), .I3(rd_addr_r_c[1]), .O(n13247));
    defparam rd_addr_r_0__bdd_4_lut_11250.LUT_INIT = 16'he4aa;
    SB_LUT4 n13247_bdd_4_lut (.I0(n13247), .I1(\REG.mem_17_6 ), .I2(\REG.mem_16_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11110));
    defparam n13247_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3882_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_21_7 ), .O(n5265));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3882_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3881_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_21_6 ), .O(n5264));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3881_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3880_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_21_5 ), .O(n5263));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3880_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3879_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_21_4 ), .O(n5262));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3879_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3878_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_21_3 ), .O(n5261));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3878_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12329_bdd_4_lut (.I0(n12329), .I1(\REG.mem_9_9 ), .I2(\REG.mem_8_9 ), 
            .I3(rd_addr_r_c[1]), .O(n11158));
    defparam n12329_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11245 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_3 ), 
            .I2(\REG.mem_51_3 ), .I3(rd_addr_r_c[1]), .O(n13241));
    defparam rd_addr_r_0__bdd_4_lut_11245.LUT_INIT = 16'he4aa;
    SB_LUT4 n12599_bdd_4_lut (.I0(n12599), .I1(n11719), .I2(n11710), .I3(rd_addr_r_c[3]), 
            .O(n11767));
    defparam n12599_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13241_bdd_4_lut (.I0(n13241), .I1(\REG.mem_49_3 ), .I2(\REG.mem_48_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11113));
    defparam n13241_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3877_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_21_2 ), .O(n5260));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3877_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3876_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_21_1 ), .O(n5259));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3876_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10712 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_0 ), 
            .I2(\REG.mem_43_0 ), .I3(rd_addr_r_c[1]), .O(n12593));
    defparam rd_addr_r_0__bdd_4_lut_10712.LUT_INIT = 16'he4aa;
    SB_LUT4 i3874_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_21_0 ), .O(n5257));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3874_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3906_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_22_15 ), .O(n5289));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3906_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3905_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_22_14 ), .O(n5288));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3905_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3904_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_22_13 ), .O(n5287));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3904_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11270 (.I0(rd_addr_r_c[1]), .I1(n11996), 
            .I2(n11997), .I3(rd_addr_r_c[2]), .O(n13235));
    defparam rd_addr_r_1__bdd_4_lut_11270.LUT_INIT = 16'he4aa;
    SB_LUT4 n12593_bdd_4_lut (.I0(n12593), .I1(\REG.mem_41_0 ), .I2(\REG.mem_40_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11335));
    defparam n12593_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13235_bdd_4_lut (.I0(n13235), .I1(n11991), .I2(n11990), .I3(rd_addr_r_c[2]), 
            .O(n13238));
    defparam n13235_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3903_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_22_12 ), .O(n5286));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3903_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3902_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_22_11 ), .O(n5285));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3902_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3901_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_22_10 ), .O(n5284));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3901_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3900_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_22_9 ), .O(n5283));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3900_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3899_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_22_8 ), .O(n5282));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3899_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3898_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_22_7 ), .O(n5281));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3898_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3897_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_22_6 ), .O(n5280));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3897_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3896_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_22_5 ), .O(n5279));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3896_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3895_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_22_4 ), .O(n5278));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3895_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3894_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_22_3 ), .O(n5277));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3894_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3893_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_22_2 ), .O(n5276));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3893_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11240 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_11 ), 
            .I2(\REG.mem_15_11 ), .I3(rd_addr_r_c[1]), .O(n13229));
    defparam rd_addr_r_0__bdd_4_lut_11240.LUT_INIT = 16'he4aa;
    SB_LUT4 i3892_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_22_1 ), .O(n5275));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3892_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13229_bdd_4_lut (.I0(n13229), .I1(\REG.mem_13_11 ), .I2(\REG.mem_12_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11632));
    defparam n13229_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3891_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_22_0 ), .O(n5274));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3891_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3946_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_24_15 ), .O(n5329));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3946_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_10622 (.I0(rd_addr_r_c[4]), .I1(n11728), 
            .I2(n11785), .I3(rd_addr_r_c[5]), .O(n12401));
    defparam rd_addr_r_4__bdd_4_lut_10622.LUT_INIT = 16'he4aa;
    SB_LUT4 i3945_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_24_14 ), .O(n5328));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3945_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3944_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_24_13 ), .O(n5327));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3944_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12401_bdd_4_lut (.I0(n12401), .I1(n11704), .I2(n11659), .I3(rd_addr_r_c[5]), 
            .O(\REG.out_raw_31__N_559 [6]));
    defparam n12401_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3943_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_24_12 ), .O(n5326));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3943_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11230 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_13 ), 
            .I2(\REG.mem_59_13 ), .I3(rd_addr_r_c[1]), .O(n13223));
    defparam rd_addr_r_0__bdd_4_lut_11230.LUT_INIT = 16'he4aa;
    SB_LUT4 i3942_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_24_11 ), .O(n5325));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3942_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10702 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_5 ), 
            .I2(\REG.mem_39_5 ), .I3(rd_addr_r_c[1]), .O(n12581));
    defparam rd_addr_r_0__bdd_4_lut_10702.LUT_INIT = 16'he4aa;
    SB_LUT4 n12581_bdd_4_lut (.I0(n12581), .I1(\REG.mem_37_5 ), .I2(\REG.mem_36_5 ), 
            .I3(rd_addr_r_c[1]), .O(n12584));
    defparam n12581_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13223_bdd_4_lut (.I0(n13223), .I1(\REG.mem_57_13 ), .I2(\REG.mem_56_13 ), 
            .I3(rd_addr_r_c[1]), .O(n13226));
    defparam n13223_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11235 (.I0(rd_addr_r_c[1]), .I1(n11240), 
            .I2(n11241), .I3(rd_addr_r_c[2]), .O(n13217));
    defparam rd_addr_r_1__bdd_4_lut_11235.LUT_INIT = 16'he4aa;
    SB_LUT4 i3941_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_24_10 ), .O(n5324));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3941_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i56_57 (.Q(\REG.mem_0_6 ), .C(FIFO_CLK_c), .D(n4933));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3940_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_24_9 ), .O(n5323));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3940_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \REG.out_buffer__i2  (.Q(\fifo_data_out[2] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n6121));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 n13217_bdd_4_lut (.I0(n13217), .I1(n11238), .I2(n11237), .I3(rd_addr_r_c[2]), 
            .O(n11262));
    defparam n13217_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \REG.out_buffer__i1  (.Q(\fifo_data_out[1] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n6118));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 i3939_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_24_8 ), .O(n5322));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3939_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3938_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_24_7 ), .O(n5321));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3938_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11225 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_1 ), 
            .I2(\REG.mem_51_1 ), .I3(rd_addr_r_c[1]), .O(n13211));
    defparam rd_addr_r_0__bdd_4_lut_11225.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10692 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_9 ), 
            .I2(\REG.mem_7_9 ), .I3(rd_addr_r_c[1]), .O(n12575));
    defparam rd_addr_r_0__bdd_4_lut_10692.LUT_INIT = 16'he4aa;
    SB_LUT4 i3937_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_24_6 ), .O(n5320));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3937_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13211_bdd_4_lut (.I0(n13211), .I1(\REG.mem_49_1 ), .I2(\REG.mem_48_1 ), 
            .I3(rd_addr_r_c[1]), .O(n13214));
    defparam n13211_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF \REG.out_buffer__i3  (.Q(\fifo_data_out[3] ), .C(SLM_CLK_c), 
           .D(n10556));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i4  (.Q(\fifo_data_out[4] ), .C(SLM_CLK_c), 
           .D(n10562));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i4_1_lut (.I0(rd_addr_r_c[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11215 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_11 ), 
            .I2(\REG.mem_19_11 ), .I3(rd_addr_r_c[1]), .O(n13205));
    defparam rd_addr_r_0__bdd_4_lut_11215.LUT_INIT = 16'he4aa;
    SB_LUT4 i4369_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_49_15 ), .O(n5752));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4369_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13205_bdd_4_lut (.I0(n13205), .I1(\REG.mem_17_11 ), .I2(\REG.mem_16_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11644));
    defparam n13205_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9545_3_lut (.I0(n12956), .I1(n12308), .I2(rd_addr_r_c[3]), 
            .I3(GND_net), .O(n11383));
    defparam i9545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4368_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_49_14 ), .O(n5751));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4368_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3936_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_24_5 ), .O(n5319));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3936_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3935_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_24_4 ), .O(n5318));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3935_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3934_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_24_3 ), .O(n5317));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3934_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3933_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_24_2 ), .O(n5316));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3933_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12575_bdd_4_lut (.I0(n12575), .I1(\REG.mem_5_9 ), .I2(\REG.mem_4_9 ), 
            .I3(rd_addr_r_c[1]), .O(n11143));
    defparam n12575_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3932_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_24_1 ), .O(n5315));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3932_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF \REG.out_buffer__i5  (.Q(\fifo_data_out[5] ), .C(SLM_CLK_c), 
           .D(n10564));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 i3924_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_24_0 ), .O(n5307));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3924_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF \REG.out_buffer__i6  (.Q(\fifo_data_out[6] ), .C(SLM_CLK_c), 
           .D(n10566));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i7  (.Q(\fifo_data_out[7] ), .C(SLM_CLK_c), 
           .D(n10568));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i8  (.Q(\fifo_data_out[8] ), .C(SLM_CLK_c), 
           .D(n10570));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i9  (.Q(\fifo_data_out[9] ), .C(SLM_CLK_c), 
           .D(n10572));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i10  (.Q(\fifo_data_out[10] ), .C(SLM_CLK_c), 
           .D(n10574));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i11  (.Q(\fifo_data_out[11] ), .C(SLM_CLK_c), 
           .D(n10576));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 i4367_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_49_13 ), .O(n5750));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4367_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3978_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_26_15 ), .O(n5361));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3978_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4366_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_49_12 ), .O(n5749));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4366_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3977_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_26_14 ), .O(n5360));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3977_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4365_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_49_11 ), .O(n5748));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4365_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11210 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_5 ), 
            .I2(\REG.mem_31_5 ), .I3(rd_addr_r_c[1]), .O(n13199));
    defparam rd_addr_r_0__bdd_4_lut_11210.LUT_INIT = 16'he4aa;
    SB_LUT4 i4364_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_49_10 ), .O(n5747));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4364_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13199_bdd_4_lut (.I0(n13199), .I1(\REG.mem_29_5 ), .I2(\REG.mem_28_5 ), 
            .I3(rd_addr_r_c[1]), .O(n13202));
    defparam n13199_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \REG.out_buffer__i0  (.Q(\fifo_data_out[0] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n6085));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 i4363_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_49_9 ), .O(n5746));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4363_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4362_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_49_8 ), .O(n5745));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4362_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11205 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_12 ), 
            .I2(\REG.mem_27_12 ), .I3(rd_addr_r_c[1]), .O(n13193));
    defparam rd_addr_r_0__bdd_4_lut_11205.LUT_INIT = 16'he4aa;
    SB_LUT4 i3976_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_26_13 ), .O(n5359));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3976_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3975_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_26_12 ), .O(n5358));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3975_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4361_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_49_7 ), .O(n5744));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4361_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13193_bdd_4_lut (.I0(n13193), .I1(\REG.mem_25_12 ), .I2(\REG.mem_24_12 ), 
            .I3(rd_addr_r_c[1]), .O(n13196));
    defparam n13193_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i6_1_lut (.I0(rd_addr_r_c[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10548 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_13 ), 
            .I2(\REG.mem_39_13 ), .I3(rd_addr_r_c[1]), .O(n12395));
    defparam rd_addr_r_0__bdd_4_lut_10548.LUT_INIT = 16'he4aa;
    SB_LUT4 i4360_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_49_6 ), .O(n5743));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4360_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4359_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_49_5 ), .O(n5742));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4359_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3974_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_26_11 ), .O(n5357));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3974_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4358_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_49_4 ), .O(n5741));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4358_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF \REG.out_buffer__i12  (.Q(\fifo_data_out[12] ), .C(SLM_CLK_c), 
           .D(n10578));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i13  (.Q(\fifo_data_out[13] ), .C(SLM_CLK_c), 
           .D(n10580));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF i59_60 (.Q(\REG.mem_0_7 ), .C(FIFO_CLK_c), .D(n4932));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4357_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_49_3 ), .O(n5740));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4357_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wp_sync2_r_6__I_0_143_i1_2_lut (.I0(wp_sync2_r[5]), .I1(wp_sync2_r[6]), 
            .I2(GND_net), .I3(GND_net), .O(wp_sync_w[5]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam wp_sync2_r_6__I_0_143_i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3973_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_26_10 ), .O(n5356));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3973_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3972_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_26_9 ), .O(n5355));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3972_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i7_1_lut (.I0(\rd_addr_r[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3971_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_26_8 ), .O(n5354));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3971_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3970_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_26_7 ), .O(n5353));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3970_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4356_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_49_2 ), .O(n5739));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4356_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3969_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_26_6 ), .O(n5352));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3969_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11200 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_15 ), 
            .I2(\REG.mem_7_15 ), .I3(rd_addr_r_c[1]), .O(n13187));
    defparam rd_addr_r_0__bdd_4_lut_11200.LUT_INIT = 16'he4aa;
    SB_LUT4 i4355_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_49_1 ), .O(n5738));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4355_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3968_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_26_5 ), .O(n5351));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3968_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF wr_addr_r__i1 (.Q(wr_addr_r[1]), .C(FIFO_CLK_c), .D(n6045));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i2 (.Q(wr_addr_r[2]), .C(FIFO_CLK_c), .D(n6044));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i3 (.Q(wr_addr_r[3]), .C(FIFO_CLK_c), .D(n6043));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i4 (.Q(wr_addr_r[4]), .C(FIFO_CLK_c), .D(n6042));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 n13187_bdd_4_lut (.I0(n13187), .I1(\REG.mem_5_15 ), .I2(\REG.mem_4_15 ), 
            .I3(rd_addr_r_c[1]), .O(n13190));
    defparam n13187_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4354_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_49_0 ), .O(n5737));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4354_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11195 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_13 ), 
            .I2(\REG.mem_35_13 ), .I3(rd_addr_r_c[1]), .O(n13181));
    defparam rd_addr_r_0__bdd_4_lut_11195.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10707 (.I0(rd_addr_r_c[2]), .I1(n11335), 
            .I2(n11947), .I3(rd_addr_r_c[3]), .O(n12551));
    defparam rd_addr_r_2__bdd_4_lut_10707.LUT_INIT = 16'he4aa;
    SB_DFF wr_addr_r__i5 (.Q(wr_addr_r[5]), .C(FIFO_CLK_c), .D(n6024));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF i6131_6132 (.Q(\REG.mem_63_15 ), .C(FIFO_CLK_c), .D(n6021));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6128_6129 (.Q(\REG.mem_63_14 ), .C(FIFO_CLK_c), .D(n6020));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6125_6126 (.Q(\REG.mem_63_13 ), .C(FIFO_CLK_c), .D(n6019));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6122_6123 (.Q(\REG.mem_63_12 ), .C(FIFO_CLK_c), .D(n6018));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i62_63 (.Q(\REG.mem_0_8 ), .C(FIFO_CLK_c), .D(n4931));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12551_bdd_4_lut (.I0(n12551), .I1(n11332), .I2(n11320), .I3(rd_addr_r_c[3]), 
            .O(n12554));
    defparam n12551_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13181_bdd_4_lut (.I0(n13181), .I1(\REG.mem_33_13 ), .I2(\REG.mem_32_13 ), 
            .I3(rd_addr_r_c[1]), .O(n13184));
    defparam n13181_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11190 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_6 ), 
            .I2(\REG.mem_27_6 ), .I3(rd_addr_r_c[1]), .O(n13175));
    defparam rd_addr_r_0__bdd_4_lut_11190.LUT_INIT = 16'he4aa;
    SB_LUT4 i3967_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_26_4 ), .O(n5350));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3967_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i6119_6120 (.Q(\REG.mem_63_11 ), .C(FIFO_CLK_c), .D(n6017));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10667 (.I0(rd_addr_r_c[2]), .I1(n11089), 
            .I2(n11104), .I3(rd_addr_r_c[3]), .O(n12545));
    defparam rd_addr_r_2__bdd_4_lut_10667.LUT_INIT = 16'he4aa;
    SB_LUT4 i3966_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_26_3 ), .O(n5349));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3966_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i6116_6117 (.Q(\REG.mem_63_10 ), .C(FIFO_CLK_c), .D(n6016));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6113_6114 (.Q(\REG.mem_63_9 ), .C(FIFO_CLK_c), .D(n6015));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6110_6111 (.Q(\REG.mem_63_8 ), .C(FIFO_CLK_c), .D(n6014));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6107_6108 (.Q(\REG.mem_63_7 ), .C(FIFO_CLK_c), .D(n6013));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6104_6105 (.Q(\REG.mem_63_6 ), .C(FIFO_CLK_c), .D(n6012));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6101_6102 (.Q(\REG.mem_63_5 ), .C(FIFO_CLK_c), .D(n6011));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6098_6099 (.Q(\REG.mem_63_4 ), .C(FIFO_CLK_c), .D(n6010));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6095_6096 (.Q(\REG.mem_63_3 ), .C(FIFO_CLK_c), .D(n6009));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6092_6093 (.Q(\REG.mem_63_2 ), .C(FIFO_CLK_c), .D(n6008));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6089_6090 (.Q(\REG.mem_63_1 ), .C(FIFO_CLK_c), .D(n6007));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6086_6087 (.Q(\REG.mem_63_0 ), .C(FIFO_CLK_c), .D(n6006));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6035_6036 (.Q(\REG.mem_62_15 ), .C(FIFO_CLK_c), .D(n6005));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6032_6033 (.Q(\REG.mem_62_14 ), .C(FIFO_CLK_c), .D(n6004));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6029_6030 (.Q(\REG.mem_62_13 ), .C(FIFO_CLK_c), .D(n6003));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6026_6027 (.Q(\REG.mem_62_12 ), .C(FIFO_CLK_c), .D(n6002));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i65_66 (.Q(\REG.mem_0_9 ), .C(FIFO_CLK_c), .D(n4930));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13175_bdd_4_lut (.I0(n13175), .I1(\REG.mem_25_6 ), .I2(\REG.mem_24_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11272));
    defparam n13175_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12395_bdd_4_lut (.I0(n12395), .I1(\REG.mem_37_13 ), .I2(\REG.mem_36_13 ), 
            .I3(rd_addr_r_c[1]), .O(n12398));
    defparam n12395_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12545_bdd_4_lut (.I0(n12545), .I1(n11086), .I2(n11080), .I3(rd_addr_r_c[3]), 
            .O(n11146));
    defparam n12545_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3965_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_26_2 ), .O(n5348));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3965_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9399_3_lut (.I0(\REG.mem_56_4 ), .I1(\REG.mem_57_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11237));
    defparam i9399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10687 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_7 ), 
            .I2(\REG.mem_19_7 ), .I3(rd_addr_r_c[1]), .O(n12539));
    defparam rd_addr_r_0__bdd_4_lut_10687.LUT_INIT = 16'he4aa;
    SB_LUT4 n12539_bdd_4_lut (.I0(n12539), .I1(\REG.mem_17_7 ), .I2(\REG.mem_16_7 ), 
            .I3(rd_addr_r_c[1]), .O(n12542));
    defparam n12539_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9400_3_lut (.I0(\REG.mem_58_4 ), .I1(\REG.mem_59_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11238));
    defparam i9400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10662 (.I0(rd_addr_r_c[2]), .I1(n11593), 
            .I2(n11614), .I3(rd_addr_r_c[3]), .O(n12533));
    defparam rd_addr_r_2__bdd_4_lut_10662.LUT_INIT = 16'he4aa;
    SB_DFF i68_69 (.Q(\REG.mem_0_10 ), .C(FIFO_CLK_c), .D(n4929));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i71_72 (.Q(\REG.mem_0_11 ), .C(FIFO_CLK_c), .D(n4928));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12533_bdd_4_lut (.I0(n12533), .I1(n11545), .I2(n11530), .I3(rd_addr_r_c[3]), 
            .O(n11785));
    defparam n12533_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i6023_6024 (.Q(\REG.mem_62_11 ), .C(FIFO_CLK_c), .D(n6001));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6020_6021 (.Q(\REG.mem_62_10 ), .C(FIFO_CLK_c), .D(n6000));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6017_6018 (.Q(\REG.mem_62_9 ), .C(FIFO_CLK_c), .D(n5999));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6014_6015 (.Q(\REG.mem_62_8 ), .C(FIFO_CLK_c), .D(n5998));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6011_6012 (.Q(\REG.mem_62_7 ), .C(FIFO_CLK_c), .D(n5997));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6008_6009 (.Q(\REG.mem_62_6 ), .C(FIFO_CLK_c), .D(n5996));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6005_6006 (.Q(\REG.mem_62_5 ), .C(FIFO_CLK_c), .D(n5995));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6002_6003 (.Q(\REG.mem_62_4 ), .C(FIFO_CLK_c), .D(n5994));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5999_6000 (.Q(\REG.mem_62_3 ), .C(FIFO_CLK_c), .D(n5993));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5996_5997 (.Q(\REG.mem_62_2 ), .C(FIFO_CLK_c), .D(n5992));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5993_5994 (.Q(\REG.mem_62_1 ), .C(FIFO_CLK_c), .D(n5991));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5990_5991 (.Q(\REG.mem_62_0 ), .C(FIFO_CLK_c), .D(n5990));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5939_5940 (.Q(\REG.mem_61_15 ), .C(FIFO_CLK_c), .D(n5986));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5936_5937 (.Q(\REG.mem_61_14 ), .C(FIFO_CLK_c), .D(n5985));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3964_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_26_1 ), .O(n5347));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3964_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10657 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_15 ), 
            .I2(\REG.mem_39_15 ), .I3(rd_addr_r_c[1]), .O(n12527));
    defparam rd_addr_r_0__bdd_4_lut_10657.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11185 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_11 ), 
            .I2(\REG.mem_23_11 ), .I3(rd_addr_r_c[1]), .O(n13169));
    defparam rd_addr_r_0__bdd_4_lut_11185.LUT_INIT = 16'he4aa;
    SB_LUT4 n12527_bdd_4_lut (.I0(n12527), .I1(\REG.mem_37_15 ), .I2(\REG.mem_36_15 ), 
            .I3(rd_addr_r_c[1]), .O(n12530));
    defparam n12527_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3963_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_26_0 ), .O(n5346));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3963_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13169_bdd_4_lut (.I0(n13169), .I1(\REG.mem_21_11 ), .I2(\REG.mem_20_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11653));
    defparam n13169_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10652 (.I0(rd_addr_r_c[2]), .I1(n11125), 
            .I2(n11128), .I3(rd_addr_r_c[3]), .O(n12521));
    defparam rd_addr_r_2__bdd_4_lut_10652.LUT_INIT = 16'he4aa;
    SB_LUT4 n12521_bdd_4_lut (.I0(n12521), .I1(n11119), .I2(n11113), .I3(rd_addr_r_c[3]), 
            .O(n11149));
    defparam n12521_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_11495 (.I0(rd_addr_r_c[4]), .I1(n11146), 
            .I2(n11149), .I3(rd_addr_r_c[5]), .O(n12515));
    defparam rd_addr_r_4__bdd_4_lut_11495.LUT_INIT = 16'he4aa;
    SB_LUT4 n12515_bdd_4_lut (.I0(n12515), .I1(n11137), .I2(n11131), .I3(rd_addr_r_c[5]), 
            .O(\REG.out_raw_31__N_559 [3]));
    defparam n12515_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i5933_5934 (.Q(\REG.mem_61_13 ), .C(FIFO_CLK_c), .D(n5984));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5930_5931 (.Q(\REG.mem_61_12 ), .C(FIFO_CLK_c), .D(n5983));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5927_5928 (.Q(\REG.mem_61_11 ), .C(FIFO_CLK_c), .D(n5982));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5924_5925 (.Q(\REG.mem_61_10 ), .C(FIFO_CLK_c), .D(n5981));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5921_5922 (.Q(\REG.mem_61_9 ), .C(FIFO_CLK_c), .D(n5980));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5918_5919 (.Q(\REG.mem_61_8 ), .C(FIFO_CLK_c), .D(n5979));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5915_5916 (.Q(\REG.mem_61_7 ), .C(FIFO_CLK_c), .D(n5978));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5912_5913 (.Q(\REG.mem_61_6 ), .C(FIFO_CLK_c), .D(n5977));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5909_5910 (.Q(\REG.mem_61_5 ), .C(FIFO_CLK_c), .D(n5976));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5906_5907 (.Q(\REG.mem_61_4 ), .C(FIFO_CLK_c), .D(n5975));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5903_5904 (.Q(\REG.mem_61_3 ), .C(FIFO_CLK_c), .D(n5974));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5900_5901 (.Q(\REG.mem_61_2 ), .C(FIFO_CLK_c), .D(n5973));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5897_5898 (.Q(\REG.mem_61_1 ), .C(FIFO_CLK_c), .D(n5972));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5894_5895 (.Q(\REG.mem_61_0 ), .C(FIFO_CLK_c), .D(n5971));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5843_5844 (.Q(\REG.mem_60_15 ), .C(FIFO_CLK_c), .D(n5969));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11180 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_11 ), 
            .I2(\REG.mem_27_11 ), .I3(rd_addr_r_c[1]), .O(n13163));
    defparam rd_addr_r_0__bdd_4_lut_11180.LUT_INIT = 16'he4aa;
    SB_LUT4 n13163_bdd_4_lut (.I0(n13163), .I1(\REG.mem_25_11 ), .I2(\REG.mem_24_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11656));
    defparam n13163_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3994_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_27_15 ), .O(n5377));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3994_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3993_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_27_14 ), .O(n5376));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3993_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10647 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_12 ), 
            .I2(\REG.mem_59_12 ), .I3(rd_addr_r_c[1]), .O(n12509));
    defparam rd_addr_r_0__bdd_4_lut_10647.LUT_INIT = 16'he4aa;
    SB_LUT4 i9403_3_lut (.I0(\REG.mem_62_4 ), .I1(\REG.mem_63_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11241));
    defparam i9403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9402_3_lut (.I0(\REG.mem_60_4 ), .I1(\REG.mem_61_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11240));
    defparam i9402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11275 (.I0(rd_addr_r_c[3]), .I1(n12878), 
            .I2(n11262), .I3(rd_addr_r_c[4]), .O(n13157));
    defparam rd_addr_r_3__bdd_4_lut_11275.LUT_INIT = 16'he4aa;
    SB_LUT4 n12509_bdd_4_lut (.I0(n12509), .I1(\REG.mem_57_12 ), .I2(\REG.mem_56_12 ), 
            .I3(rd_addr_r_c[1]), .O(n12512));
    defparam n12509_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3992_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_27_13 ), .O(n5375));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3992_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9821_3_lut (.I0(n13142), .I1(n13148), .I2(rd_addr_r_c[3]), 
            .I3(GND_net), .O(n11659));
    defparam i9821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13157_bdd_4_lut (.I0(n13157), .I1(n11259), .I2(n12872), .I3(rd_addr_r_c[4]), 
            .O(n13160));
    defparam n13157_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i5840_5841 (.Q(\REG.mem_60_14 ), .C(FIFO_CLK_c), .D(n5968));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10152_3_lut (.I0(\REG.mem_40_14 ), .I1(\REG.mem_41_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11990));
    defparam i10152_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5837_5838 (.Q(\REG.mem_60_13 ), .C(FIFO_CLK_c), .D(n5967));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5834_5835 (.Q(\REG.mem_60_12 ), .C(FIFO_CLK_c), .D(n5966));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5831_5832 (.Q(\REG.mem_60_11 ), .C(FIFO_CLK_c), .D(n5965));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5828_5829 (.Q(\REG.mem_60_10 ), .C(FIFO_CLK_c), .D(n5964));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5825_5826 (.Q(\REG.mem_60_9 ), .C(FIFO_CLK_c), .D(n5963));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5822_5823 (.Q(\REG.mem_60_8 ), .C(FIFO_CLK_c), .D(n5962));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5819_5820 (.Q(\REG.mem_60_7 ), .C(FIFO_CLK_c), .D(n5961));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5816_5817 (.Q(\REG.mem_60_6 ), .C(FIFO_CLK_c), .D(n5960));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5813_5814 (.Q(\REG.mem_60_5 ), .C(FIFO_CLK_c), .D(n5959));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5810_5811 (.Q(\REG.mem_60_4 ), .C(FIFO_CLK_c), .D(n5958));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5807_5808 (.Q(\REG.mem_60_3 ), .C(FIFO_CLK_c), .D(n5957));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5804_5805 (.Q(\REG.mem_60_2 ), .C(FIFO_CLK_c), .D(n5956));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5801_5802 (.Q(\REG.mem_60_1 ), .C(FIFO_CLK_c), .D(n5955));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5798_5799 (.Q(\REG.mem_60_0 ), .C(FIFO_CLK_c), .D(n5954));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync1_r__i1 (.Q(rp_sync1_r[1]), .C(FIFO_CLK_c), .D(n5953));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_LUT4 i10153_3_lut (.I0(\REG.mem_42_14 ), .I1(\REG.mem_43_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11991));
    defparam i10153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10159_3_lut (.I0(\REG.mem_46_14 ), .I1(\REG.mem_47_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11997));
    defparam i10159_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF rp_sync1_r__i2 (.Q(rp_sync1_r[2]), .C(FIFO_CLK_c), .D(n5952));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i3 (.Q(rp_sync1_r[3]), .C(FIFO_CLK_c), .D(n5951));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i4 (.Q(rp_sync1_r[4]), .C(FIFO_CLK_c), .D(n5950));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i5 (.Q(rp_sync1_r[5]), .C(FIFO_CLK_c), .D(n5949));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i6 (.Q(rp_sync1_r[6]), .C(FIFO_CLK_c), .D(n5948));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i1 (.Q(rp_sync2_r[1]), .C(FIFO_CLK_c), .D(n5947));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i2 (.Q(rp_sync2_r[2]), .C(FIFO_CLK_c), .D(n5946));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i3 (.Q(rp_sync2_r[3]), .C(FIFO_CLK_c), .D(n5945));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF i5747_5748 (.Q(\REG.mem_59_15 ), .C(FIFO_CLK_c), .D(n5944));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5744_5745 (.Q(\REG.mem_59_14 ), .C(FIFO_CLK_c), .D(n5943));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5741_5742 (.Q(\REG.mem_59_13 ), .C(FIFO_CLK_c), .D(n5942));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5738_5739 (.Q(\REG.mem_59_12 ), .C(FIFO_CLK_c), .D(n5941));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5735_5736 (.Q(\REG.mem_59_11 ), .C(FIFO_CLK_c), .D(n5940));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5732_5733 (.Q(\REG.mem_59_10 ), .C(FIFO_CLK_c), .D(n5939));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5729_5730 (.Q(\REG.mem_59_9 ), .C(FIFO_CLK_c), .D(n5938));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5726_5727 (.Q(\REG.mem_59_8 ), .C(FIFO_CLK_c), .D(n5937));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10632 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_9 ), 
            .I2(\REG.mem_55_9 ), .I3(rd_addr_r_c[1]), .O(n12503));
    defparam rd_addr_r_0__bdd_4_lut_10632.LUT_INIT = 16'he4aa;
    SB_LUT4 i3991_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_27_12 ), .O(n5374));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3991_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12503_bdd_4_lut (.I0(n12503), .I1(\REG.mem_53_9 ), .I2(\REG.mem_52_9 ), 
            .I3(rd_addr_r_c[1]), .O(n12506));
    defparam n12503_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10158_3_lut (.I0(\REG.mem_44_14 ), .I1(\REG.mem_45_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11996));
    defparam i10158_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5723_5724 (.Q(\REG.mem_59_7 ), .C(FIFO_CLK_c), .D(n5936));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5720_5721 (.Q(\REG.mem_59_6 ), .C(FIFO_CLK_c), .D(n5935));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11175 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_7 ), 
            .I2(\REG.mem_11_7 ), .I3(rd_addr_r_c[1]), .O(n13151));
    defparam rd_addr_r_0__bdd_4_lut_11175.LUT_INIT = 16'he4aa;
    SB_DFF i5717_5718 (.Q(\REG.mem_59_5 ), .C(FIFO_CLK_c), .D(n5934));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5714_5715 (.Q(\REG.mem_59_4 ), .C(FIFO_CLK_c), .D(n5933));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5711_5712 (.Q(\REG.mem_59_3 ), .C(FIFO_CLK_c), .D(n5932));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5708_5709 (.Q(\REG.mem_59_2 ), .C(FIFO_CLK_c), .D(n5931));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5705_5706 (.Q(\REG.mem_59_1 ), .C(FIFO_CLK_c), .D(n5930));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5702_5703 (.Q(\REG.mem_59_0 ), .C(FIFO_CLK_c), .D(n5929));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync2_r__i4 (.Q(rp_sync2_r[4]), .C(FIFO_CLK_c), .D(n5928));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i5 (.Q(rp_sync2_r[5]), .C(FIFO_CLK_c), .D(n5927));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i6 (.Q(rp_sync2_r[6]), .C(FIFO_CLK_c), .D(n5926));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rd_addr_r__i1 (.Q(rd_addr_r_c[1]), .C(SLM_CLK_c), .D(n5925));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i2 (.Q(rd_addr_r_c[2]), .C(SLM_CLK_c), .D(n5924));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i3 (.Q(rd_addr_r_c[3]), .C(SLM_CLK_c), .D(n5923));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i4 (.Q(rd_addr_r_c[4]), .C(SLM_CLK_c), .D(n5922));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i5 (.Q(rd_addr_r_c[5]), .C(SLM_CLK_c), .D(n5921));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i6 (.Q(\rd_addr_r[6] ), .C(SLM_CLK_c), .D(n5920));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF i5651_5652 (.Q(\REG.mem_58_15 ), .C(FIFO_CLK_c), .D(n5919));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13151_bdd_4_lut (.I0(n13151), .I1(\REG.mem_9_7 ), .I2(\REG.mem_8_7 ), 
            .I3(rd_addr_r_c[1]), .O(n13154));
    defparam n13151_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i5648_5649 (.Q(\REG.mem_58_14 ), .C(FIFO_CLK_c), .D(n5918));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i74_75 (.Q(\REG.mem_0_12 ), .C(FIFO_CLK_c), .D(n4927));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_4__bdd_4_lut_10637 (.I0(rd_addr_r_c[4]), .I1(n11764), 
            .I2(n11767), .I3(rd_addr_r_c[5]), .O(n12497));
    defparam rd_addr_r_4__bdd_4_lut_10637.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11220 (.I0(rd_addr_r_c[1]), .I1(n11093), 
            .I2(n11094), .I3(rd_addr_r_c[2]), .O(n13145));
    defparam rd_addr_r_1__bdd_4_lut_11220.LUT_INIT = 16'he4aa;
    SB_LUT4 i3990_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_27_11 ), .O(n5373));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3990_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i5645_5646 (.Q(\REG.mem_58_13 ), .C(FIFO_CLK_c), .D(n5917));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5642_5643 (.Q(\REG.mem_58_12 ), .C(FIFO_CLK_c), .D(n5916));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9378_3_lut (.I0(\REG.mem_40_4 ), .I1(\REG.mem_41_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11216));
    defparam i9378_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5639_5640 (.Q(\REG.mem_58_11 ), .C(FIFO_CLK_c), .D(n5915));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5636_5637 (.Q(\REG.mem_58_10 ), .C(FIFO_CLK_c), .D(n5914));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5633_5634 (.Q(\REG.mem_58_9 ), .C(FIFO_CLK_c), .D(n5913));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5630_5631 (.Q(\REG.mem_58_8 ), .C(FIFO_CLK_c), .D(n5912));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5627_5628 (.Q(\REG.mem_58_7 ), .C(FIFO_CLK_c), .D(n5911));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5624_5625 (.Q(\REG.mem_58_6 ), .C(FIFO_CLK_c), .D(n5910));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5621_5622 (.Q(\REG.mem_58_5 ), .C(FIFO_CLK_c), .D(n5909));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5618_5619 (.Q(\REG.mem_58_4 ), .C(FIFO_CLK_c), .D(n5908));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5615_5616 (.Q(\REG.mem_58_3 ), .C(FIFO_CLK_c), .D(n5907));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5612_5613 (.Q(\REG.mem_58_2 ), .C(FIFO_CLK_c), .D(n5906));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5609_5610 (.Q(\REG.mem_58_1 ), .C(FIFO_CLK_c), .D(n5905));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5606_5607 (.Q(\REG.mem_58_0 ), .C(FIFO_CLK_c), .D(n5904));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12497_bdd_4_lut (.I0(n12497), .I1(n11755), .I2(n11743), .I3(rd_addr_r_c[5]), 
            .O(\REG.out_raw_31__N_559 [11]));
    defparam n12497_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9379_3_lut (.I0(\REG.mem_42_4 ), .I1(\REG.mem_43_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11217));
    defparam i9379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13145_bdd_4_lut (.I0(n13145), .I1(n11001), .I2(n11000), .I3(rd_addr_r_c[2]), 
            .O(n13148));
    defparam n13145_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9382_3_lut (.I0(\REG.mem_46_4 ), .I1(\REG.mem_47_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11220));
    defparam i9382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9381_3_lut (.I0(\REG.mem_44_4 ), .I1(\REG.mem_45_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11219));
    defparam i9381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3989_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_27_10 ), .O(n5372));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3989_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9166_3_lut (.I0(n12686), .I1(n12296), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11004));
    defparam i9166_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5555_5556 (.Q(\REG.mem_57_15 ), .C(FIFO_CLK_c), .D(n5901));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5552_5553 (.Q(\REG.mem_57_14 ), .C(FIFO_CLK_c), .D(n5900));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5549_5550 (.Q(\REG.mem_57_13 ), .C(FIFO_CLK_c), .D(n5899));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5546_5547 (.Q(\REG.mem_57_12 ), .C(FIFO_CLK_c), .D(n5898));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5543_5544 (.Q(\REG.mem_57_11 ), .C(FIFO_CLK_c), .D(n5897));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5540_5541 (.Q(\REG.mem_57_10 ), .C(FIFO_CLK_c), .D(n5896));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5537_5538 (.Q(\REG.mem_57_9 ), .C(FIFO_CLK_c), .D(n5895));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5534_5535 (.Q(\REG.mem_57_8 ), .C(FIFO_CLK_c), .D(n5894));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5531_5532 (.Q(\REG.mem_57_7 ), .C(FIFO_CLK_c), .D(n5893));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5528_5529 (.Q(\REG.mem_57_6 ), .C(FIFO_CLK_c), .D(n5892));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5525_5526 (.Q(\REG.mem_57_5 ), .C(FIFO_CLK_c), .D(n5891));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5522_5523 (.Q(\REG.mem_57_4 ), .C(FIFO_CLK_c), .D(n5890));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5519_5520 (.Q(\REG.mem_57_3 ), .C(FIFO_CLK_c), .D(n5889));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5516_5517 (.Q(\REG.mem_57_2 ), .C(FIFO_CLK_c), .D(n5888));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5513_5514 (.Q(\REG.mem_57_1 ), .C(FIFO_CLK_c), .D(n5887));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut (.I0(rd_addr_r[0]), .I1(\REG.mem_18_1 ), 
            .I2(\REG.mem_19_1 ), .I3(rd_addr_r_c[1]), .O(n13859));
    defparam rd_addr_r_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n13859_bdd_4_lut (.I0(n13859), .I1(\REG.mem_17_1 ), .I2(\REG.mem_16_1 ), 
            .I3(rd_addr_r_c[1]), .O(n11389));
    defparam n13859_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3988_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_27_9 ), .O(n5371));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3988_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11160 (.I0(rd_addr_r_c[1]), .I1(n12023), 
            .I2(n12024), .I3(rd_addr_r_c[2]), .O(n13139));
    defparam rd_addr_r_1__bdd_4_lut_11160.LUT_INIT = 16'he4aa;
    SB_DFF i5510_5511 (.Q(\REG.mem_57_0 ), .C(FIFO_CLK_c), .D(n5885));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3987_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_27_8 ), .O(n5370));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3987_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i5459_5460 (.Q(\REG.mem_56_15 ), .C(FIFO_CLK_c), .D(n5884));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5456_5457 (.Q(\REG.mem_56_14 ), .C(FIFO_CLK_c), .D(n5883));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5453_5454 (.Q(\REG.mem_56_13 ), .C(FIFO_CLK_c), .D(n5882));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5450_5451 (.Q(\REG.mem_56_12 ), .C(FIFO_CLK_c), .D(n5881));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5447_5448 (.Q(\REG.mem_56_11 ), .C(FIFO_CLK_c), .D(n5880));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5444_5445 (.Q(\REG.mem_56_10 ), .C(FIFO_CLK_c), .D(n5879));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5441_5442 (.Q(\REG.mem_56_9 ), .C(FIFO_CLK_c), .D(n5878));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5438_5439 (.Q(\REG.mem_56_8 ), .C(FIFO_CLK_c), .D(n5877));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5435_5436 (.Q(\REG.mem_56_7 ), .C(FIFO_CLK_c), .D(n5876));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5432_5433 (.Q(\REG.mem_56_6 ), .C(FIFO_CLK_c), .D(n5875));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5429_5430 (.Q(\REG.mem_56_5 ), .C(FIFO_CLK_c), .D(n5874));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5426_5427 (.Q(\REG.mem_56_4 ), .C(FIFO_CLK_c), .D(n5873));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5423_5424 (.Q(\REG.mem_56_3 ), .C(FIFO_CLK_c), .D(n5872));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5420_5421 (.Q(\REG.mem_56_2 ), .C(FIFO_CLK_c), .D(n5871));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5417_5418 (.Q(\REG.mem_56_1 ), .C(FIFO_CLK_c), .D(n5870));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9798_3_lut (.I0(\REG.mem_32_8 ), .I1(\REG.mem_33_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11636));
    defparam i9798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9799_3_lut (.I0(\REG.mem_34_8 ), .I1(\REG.mem_35_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11637));
    defparam i9799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13139_bdd_4_lut (.I0(n13139), .I1(n12012), .I2(n12011), .I3(rd_addr_r_c[2]), 
            .O(n13142));
    defparam n13139_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9844_3_lut (.I0(\REG.mem_38_8 ), .I1(\REG.mem_39_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11682));
    defparam i9844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11755 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_14 ), 
            .I2(\REG.mem_59_14 ), .I3(rd_addr_r_c[1]), .O(n13853));
    defparam rd_addr_r_0__bdd_4_lut_11755.LUT_INIT = 16'he4aa;
    SB_LUT4 i9843_3_lut (.I0(\REG.mem_36_8 ), .I1(\REG.mem_37_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11681));
    defparam i9843_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5414_5415 (.Q(\REG.mem_56_0 ), .C(FIFO_CLK_c), .D(n5865));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wp_sync1_r__i1 (.Q(wp_sync1_r[1]), .C(SLM_CLK_c), .D(n5864));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i2 (.Q(wp_sync1_r[2]), .C(SLM_CLK_c), .D(n5863));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i3 (.Q(wp_sync1_r[3]), .C(SLM_CLK_c), .D(n5862));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i4 (.Q(wp_sync1_r[4]), .C(SLM_CLK_c), .D(n5861));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i5 (.Q(wp_sync1_r[5]), .C(SLM_CLK_c), .D(n5860));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i6 (.Q(wp_sync1_r[6]), .C(SLM_CLK_c), .D(n5859));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF i5363_5364 (.Q(\REG.mem_55_15 ), .C(FIFO_CLK_c), .D(n5858));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5360_5361 (.Q(\REG.mem_55_14 ), .C(FIFO_CLK_c), .D(n5857));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5357_5358 (.Q(\REG.mem_55_13 ), .C(FIFO_CLK_c), .D(n5856));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5354_5355 (.Q(\REG.mem_55_12 ), .C(FIFO_CLK_c), .D(n5855));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5351_5352 (.Q(\REG.mem_55_11 ), .C(FIFO_CLK_c), .D(n5854));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5348_5349 (.Q(\REG.mem_55_10 ), .C(FIFO_CLK_c), .D(n5853));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY wr_addr_r_6__I_0_141_7 (.CI(n10137), .I0(wr_addr_r[5]), .I1(GND_net), 
            .CO(n10138));
    SB_LUT4 wr_addr_r_6__I_0_141_6_lut (.I0(GND_net), .I1(wr_addr_r[4]), 
            .I2(GND_net), .I3(n10136), .O(wr_addr_p1_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_141_6 (.CI(n10136), .I0(wr_addr_r[4]), .I1(GND_net), 
            .CO(n10137));
    SB_LUT4 wr_addr_r_6__I_0_141_5_lut (.I0(GND_net), .I1(wr_addr_r[3]), 
            .I2(GND_net), .I3(n10135), .O(wr_addr_p1_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_141_5 (.CI(n10135), .I0(wr_addr_r[3]), .I1(GND_net), 
            .CO(n10136));
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_3 (.CI(n10090), .I0(wp_sync_w[1]), 
            .I1(n1[1]), .CO(n10091));
    SB_LUT4 wr_addr_r_6__I_0_141_4_lut (.I0(GND_net), .I1(wr_addr_r[2]), 
            .I2(GND_net), .I3(n10134), .O(wr_addr_p1_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_2_lut (.I0(GND_net), .I1(wp_sync_w[0]), 
            .I2(n1[0]), .I3(VCC_net), .O(\rd_sig_diff0_w[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_141_4 (.CI(n10134), .I0(wr_addr_r[2]), .I1(GND_net), 
            .CO(n10135));
    SB_DFF i5345_5346 (.Q(\REG.mem_55_9 ), .C(FIFO_CLK_c), .D(n5852));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5342_5343 (.Q(\REG.mem_55_8 ), .C(FIFO_CLK_c), .D(n5851));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5339_5340 (.Q(\REG.mem_55_7 ), .C(FIFO_CLK_c), .D(n5850));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5336_5337 (.Q(\REG.mem_55_6 ), .C(FIFO_CLK_c), .D(n5849));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5333_5334 (.Q(\REG.mem_55_5 ), .C(FIFO_CLK_c), .D(n5848));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5330_5331 (.Q(\REG.mem_55_4 ), .C(FIFO_CLK_c), .D(n5847));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5327_5328 (.Q(\REG.mem_55_3 ), .C(FIFO_CLK_c), .D(n5846));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5324_5325 (.Q(\REG.mem_55_2 ), .C(FIFO_CLK_c), .D(n5845));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5321_5322 (.Q(\REG.mem_55_1 ), .C(FIFO_CLK_c), .D(n5844));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5318_5319 (.Q(\REG.mem_55_0 ), .C(FIFO_CLK_c), .D(n5843));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wp_sync2_r__i1 (.Q(wp_sync2_r[1]), .C(SLM_CLK_c), .D(n5842));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i2 (.Q(wp_sync2_r[2]), .C(SLM_CLK_c), .D(n5841));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i3 (.Q(wp_sync2_r[3]), .C(SLM_CLK_c), .D(n5839));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i4 (.Q(wp_sync2_r[4]), .C(SLM_CLK_c), .D(n5838));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i5 (.Q(wp_sync2_r[5]), .C(SLM_CLK_c), .D(n5837));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_LUT4 wr_addr_r_6__I_0_141_3_lut (.I0(GND_net), .I1(wr_addr_r[1]), 
            .I2(GND_net), .I3(n10133), .O(wr_addr_p1_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_r_6__I_0_151_8_lut (.I0(GND_net), .I1(\rd_addr_r[6] ), 
            .I2(GND_net), .I3(n10144), .O(rd_addr_p1_w[6])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_141_3 (.CI(n10133), .I0(wr_addr_r[1]), .I1(GND_net), 
            .CO(n10134));
    SB_LUT4 wr_addr_r_6__I_0_141_2_lut (.I0(GND_net), .I1(wr_addr_r[0]), 
            .I2(GND_net), .I3(VCC_net), .O(wr_addr_p1_w[0])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_r_6__I_0_151_7_lut (.I0(GND_net), .I1(rd_addr_r_c[5]), 
            .I2(GND_net), .I3(n10143), .O(rd_addr_p1_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_141_2 (.CI(VCC_net), .I0(wr_addr_r[0]), .I1(GND_net), 
            .CO(n10133));
    SB_LUT4 i9855_3_lut (.I0(\REG.mem_16_15 ), .I1(\REG.mem_17_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11693));
    defparam i9855_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rd_addr_r_6__I_0_151_7 (.CI(n10143), .I0(rd_addr_r_c[5]), .I1(GND_net), 
            .CO(n10144));
    SB_LUT4 i9856_3_lut (.I0(\REG.mem_18_15 ), .I1(\REG.mem_19_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11694));
    defparam i9856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_add_2_8_lut (.I0(n10979), .I1(wr_grey_sync_r[6]), 
            .I2(n1_adj_45[6]), .I3(n10101), .O(\afull_flag_impl.af_flag_nxt_w )) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i9877_3_lut (.I0(\REG.mem_22_15 ), .I1(\REG.mem_23_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11715));
    defparam i9877_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF wp_sync2_r__i6 (.Q(wp_sync2_r[6]), .C(SLM_CLK_c), .D(n5836));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF i5267_5268 (.Q(\REG.mem_54_15 ), .C(FIFO_CLK_c), .D(n5835));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5264_5265 (.Q(\REG.mem_54_14 ), .C(FIFO_CLK_c), .D(n5834));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5261_5262 (.Q(\REG.mem_54_13 ), .C(FIFO_CLK_c), .D(n5833));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5258_5259 (.Q(\REG.mem_54_12 ), .C(FIFO_CLK_c), .D(n5832));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5255_5256 (.Q(\REG.mem_54_11 ), .C(FIFO_CLK_c), .D(n5831));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5252_5253 (.Q(\REG.mem_54_10 ), .C(FIFO_CLK_c), .D(n5830));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5249_5250 (.Q(\REG.mem_54_9 ), .C(FIFO_CLK_c), .D(n5829));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5246_5247 (.Q(\REG.mem_54_8 ), .C(FIFO_CLK_c), .D(n5828));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5243_5244 (.Q(\REG.mem_54_7 ), .C(FIFO_CLK_c), .D(n5827));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5240_5241 (.Q(\REG.mem_54_6 ), .C(FIFO_CLK_c), .D(n5826));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5237_5238 (.Q(\REG.mem_54_5 ), .C(FIFO_CLK_c), .D(n5825));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5234_5235 (.Q(\REG.mem_54_4 ), .C(FIFO_CLK_c), .D(n5824));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5231_5232 (.Q(\REG.mem_54_3 ), .C(FIFO_CLK_c), .D(n5823));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5228_5229 (.Q(\REG.mem_54_2 ), .C(FIFO_CLK_c), .D(n5822));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5225_5226 (.Q(\REG.mem_54_1 ), .C(FIFO_CLK_c), .D(n5821));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9876_3_lut (.I0(\REG.mem_20_15 ), .I1(\REG.mem_21_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11714));
    defparam i9876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_add_2_7_lut (.I0(n10951), .I1(wr_addr_r[5]), 
            .I2(rp_sync_w[5]), .I3(n10100), .O(n10979)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY wr_addr_r_6__I_0_add_2_7 (.CI(n10100), .I0(wr_addr_r[5]), .I1(rp_sync_w[5]), 
            .CO(n10101));
    SB_LUT4 rd_addr_r_6__I_0_151_6_lut (.I0(GND_net), .I1(rd_addr_r_c[4]), 
            .I2(GND_net), .I3(n10142), .O(rd_addr_p1_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wr_addr_r_6__I_0_add_2_6_lut (.I0(n2_adj_22), .I1(wr_addr_r[4]), 
            .I2(rp_sync_w[4]), .I3(n10099), .O(n10925)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_6_lut.LUT_INIT = 16'hebbe;
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_2 (.CI(VCC_net), .I0(wp_sync_w[0]), 
            .I1(n1[0]), .CO(n10090));
    SB_CARRY wr_addr_r_6__I_0_add_2_6 (.CI(n10099), .I0(wr_addr_r[4]), .I1(rp_sync_w[4]), 
            .CO(n10100));
    SB_LUT4 i9354_3_lut (.I0(\REG.mem_24_4 ), .I1(\REG.mem_25_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11192));
    defparam i9354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_add_2_5_lut (.I0(GND_net), .I1(wr_addr_r[3]), 
            .I2(rp_sync_w[3]), .I3(n10098), .O(wr_sig_diff0_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_add_2_5 (.CI(n10098), .I0(wr_addr_r[3]), .I1(rp_sync_w[3]), 
            .CO(n10099));
    SB_LUT4 i9355_3_lut (.I0(\REG.mem_26_4 ), .I1(\REG.mem_27_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11193));
    defparam i9355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10068_3_lut (.I0(\REG.mem_32_2 ), .I1(\REG.mem_33_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11906));
    defparam i10068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10069_3_lut (.I0(\REG.mem_34_2 ), .I1(\REG.mem_35_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11907));
    defparam i10069_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rd_addr_r_6__I_0_151_6 (.CI(n10142), .I0(rd_addr_r_c[4]), .I1(GND_net), 
            .CO(n10143));
    SB_LUT4 i9361_3_lut (.I0(\REG.mem_30_4 ), .I1(\REG.mem_31_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11199));
    defparam i9361_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5222_5223 (.Q(\REG.mem_54_0 ), .C(FIFO_CLK_c), .D(n5820));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5171_5172 (.Q(\REG.mem_53_15 ), .C(FIFO_CLK_c), .D(n5819));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5168_5169 (.Q(\REG.mem_53_14 ), .C(FIFO_CLK_c), .D(n5818));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5165_5166 (.Q(\REG.mem_53_13 ), .C(FIFO_CLK_c), .D(n5817));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5162_5163 (.Q(\REG.mem_53_12 ), .C(FIFO_CLK_c), .D(n5816));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5159_5160 (.Q(\REG.mem_53_11 ), .C(FIFO_CLK_c), .D(n5815));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5156_5157 (.Q(\REG.mem_53_10 ), .C(FIFO_CLK_c), .D(n5814));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5153_5154 (.Q(\REG.mem_53_9 ), .C(FIFO_CLK_c), .D(n5813));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5150_5151 (.Q(\REG.mem_53_8 ), .C(FIFO_CLK_c), .D(n5812));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5147_5148 (.Q(\REG.mem_53_7 ), .C(FIFO_CLK_c), .D(n5811));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5144_5145 (.Q(\REG.mem_53_6 ), .C(FIFO_CLK_c), .D(n5810));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5141_5142 (.Q(\REG.mem_53_5 ), .C(FIFO_CLK_c), .D(n5809));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5138_5139 (.Q(\REG.mem_53_4 ), .C(FIFO_CLK_c), .D(n5808));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5135_5136 (.Q(\REG.mem_53_3 ), .C(FIFO_CLK_c), .D(n5807));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5132_5133 (.Q(\REG.mem_53_2 ), .C(FIFO_CLK_c), .D(n5806));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5129_5130 (.Q(\REG.mem_53_1 ), .C(FIFO_CLK_c), .D(n5805));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9360_3_lut (.I0(\REG.mem_28_4 ), .I1(\REG.mem_29_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11198));
    defparam i9360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10072_3_lut (.I0(\REG.mem_38_2 ), .I1(\REG.mem_39_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11910));
    defparam i10072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_6__I_0_151_5_lut (.I0(GND_net), .I1(rd_addr_r_c[3]), 
            .I2(GND_net), .I3(n10141), .O(rd_addr_p1_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10071_3_lut (.I0(\REG.mem_36_2 ), .I1(\REG.mem_37_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11909));
    defparam i10071_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rd_addr_r_6__I_0_151_5 (.CI(n10141), .I0(rd_addr_r_c[3]), .I1(GND_net), 
            .CO(n10142));
    SB_DFF i5126_5127 (.Q(\REG.mem_53_0 ), .C(FIFO_CLK_c), .D(n5804));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5075_5076 (.Q(\REG.mem_52_15 ), .C(FIFO_CLK_c), .D(n5803));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5072_5073 (.Q(\REG.mem_52_14 ), .C(FIFO_CLK_c), .D(n5802));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5069_5070 (.Q(\REG.mem_52_13 ), .C(FIFO_CLK_c), .D(n5801));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5066_5067 (.Q(\REG.mem_52_12 ), .C(FIFO_CLK_c), .D(n5800));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5063_5064 (.Q(\REG.mem_52_11 ), .C(FIFO_CLK_c), .D(n5799));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5060_5061 (.Q(\REG.mem_52_10 ), .C(FIFO_CLK_c), .D(n5798));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5057_5058 (.Q(\REG.mem_52_9 ), .C(FIFO_CLK_c), .D(n5797));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5054_5055 (.Q(\REG.mem_52_8 ), .C(FIFO_CLK_c), .D(n5796));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5051_5052 (.Q(\REG.mem_52_7 ), .C(FIFO_CLK_c), .D(n5795));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5048_5049 (.Q(\REG.mem_52_6 ), .C(FIFO_CLK_c), .D(n5794));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5045_5046 (.Q(\REG.mem_52_5 ), .C(FIFO_CLK_c), .D(n5793));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5042_5043 (.Q(\REG.mem_52_4 ), .C(FIFO_CLK_c), .D(n5792));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5039_5040 (.Q(\REG.mem_52_3 ), .C(FIFO_CLK_c), .D(n5791));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5036_5037 (.Q(\REG.mem_52_2 ), .C(FIFO_CLK_c), .D(n5790));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5033_5034 (.Q(\REG.mem_52_1 ), .C(FIFO_CLK_c), .D(n5789));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11165 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_15 ), 
            .I2(\REG.mem_11_15 ), .I3(rd_addr_r_c[1]), .O(n13133));
    defparam rd_addr_r_0__bdd_4_lut_11165.LUT_INIT = 16'he4aa;
    SB_LUT4 i10104_3_lut (.I0(\REG.mem_48_2 ), .I1(\REG.mem_49_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11942));
    defparam i10104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3986_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_27_7 ), .O(n5369));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3986_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10105_3_lut (.I0(\REG.mem_50_2 ), .I1(\REG.mem_51_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11943));
    defparam i10105_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13853_bdd_4_lut (.I0(n13853), .I1(\REG.mem_57_14 ), .I2(\REG.mem_56_14 ), 
            .I3(rd_addr_r_c[1]), .O(n10993));
    defparam n13853_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10111_3_lut (.I0(\REG.mem_54_2 ), .I1(\REG.mem_55_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11949));
    defparam i10111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_add_2_4_lut (.I0(GND_net), .I1(wr_addr_r[2]), 
            .I2(rp_sync_w[2]), .I3(n10097), .O(wr_sig_diff0_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF i5030_5031 (.Q(\REG.mem_52_0 ), .C(FIFO_CLK_c), .D(n5788));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY wr_addr_r_6__I_0_add_2_4 (.CI(n10097), .I0(wr_addr_r[2]), .I1(rp_sync_w[2]), 
            .CO(n10098));
    SB_DFF i4979_4980 (.Q(\REG.mem_51_15 ), .C(FIFO_CLK_c), .D(n5787));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4976_4977 (.Q(\REG.mem_51_14 ), .C(FIFO_CLK_c), .D(n5786));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4973_4974 (.Q(\REG.mem_51_13 ), .C(FIFO_CLK_c), .D(n5785));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4970_4971 (.Q(\REG.mem_51_12 ), .C(FIFO_CLK_c), .D(n5784));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4967_4968 (.Q(\REG.mem_51_11 ), .C(FIFO_CLK_c), .D(n5783));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4964_4965 (.Q(\REG.mem_51_10 ), .C(FIFO_CLK_c), .D(n5782));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4961_4962 (.Q(\REG.mem_51_9 ), .C(FIFO_CLK_c), .D(n5781));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4958_4959 (.Q(\REG.mem_51_8 ), .C(FIFO_CLK_c), .D(n5780));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4955_4956 (.Q(\REG.mem_51_7 ), .C(FIFO_CLK_c), .D(n5779));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4952_4953 (.Q(\REG.mem_51_6 ), .C(FIFO_CLK_c), .D(n5778));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4949_4950 (.Q(\REG.mem_51_5 ), .C(FIFO_CLK_c), .D(n5777));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4946_4947 (.Q(\REG.mem_51_4 ), .C(FIFO_CLK_c), .D(n5776));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4943_4944 (.Q(\REG.mem_51_3 ), .C(FIFO_CLK_c), .D(n5775));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4940_4941 (.Q(\REG.mem_51_2 ), .C(FIFO_CLK_c), .D(n5774));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4937_4938 (.Q(\REG.mem_51_1 ), .C(FIFO_CLK_c), .D(n5773));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10110_3_lut (.I0(\REG.mem_52_2 ), .I1(\REG.mem_53_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11948));
    defparam i10110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_add_2_3_lut (.I0(GND_net), .I1(wr_addr_r[1]), 
            .I2(rp_sync_w[1]), .I3(n10096), .O(wr_sig_diff0_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_add_2_3 (.CI(n10096), .I0(wr_addr_r[1]), .I1(rp_sync_w[1]), 
            .CO(n10097));
    SB_LUT4 i9330_3_lut (.I0(\REG.mem_8_4 ), .I1(\REG.mem_9_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11168));
    defparam i9330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9331_3_lut (.I0(\REG.mem_10_4 ), .I1(\REG.mem_11_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11169));
    defparam i9331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_6__I_0_151_4_lut (.I0(GND_net), .I1(rd_addr_r_c[2]), 
            .I2(GND_net), .I3(n10140), .O(rd_addr_p1_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wr_addr_r_6__I_0_add_2_2_lut (.I0(GND_net), .I1(wr_addr_r[0]), 
            .I2(rp_sync_w[0]), .I3(VCC_net), .O(wr_sig_diff0_w[0])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF i4934_4935 (.Q(\REG.mem_51_0 ), .C(FIFO_CLK_c), .D(n5772));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4883_4884 (.Q(\REG.mem_50_15 ), .C(FIFO_CLK_c), .D(n5771));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4880_4881 (.Q(\REG.mem_50_14 ), .C(FIFO_CLK_c), .D(n5770));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4877_4878 (.Q(\REG.mem_50_13 ), .C(FIFO_CLK_c), .D(n5769));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4874_4875 (.Q(\REG.mem_50_12 ), .C(FIFO_CLK_c), .D(n5768));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4871_4872 (.Q(\REG.mem_50_11 ), .C(FIFO_CLK_c), .D(n5767));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4868_4869 (.Q(\REG.mem_50_10 ), .C(FIFO_CLK_c), .D(n5766));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4865_4866 (.Q(\REG.mem_50_9 ), .C(FIFO_CLK_c), .D(n5765));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4862_4863 (.Q(\REG.mem_50_8 ), .C(FIFO_CLK_c), .D(n5764));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4859_4860 (.Q(\REG.mem_50_7 ), .C(FIFO_CLK_c), .D(n5763));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4856_4857 (.Q(\REG.mem_50_6 ), .C(FIFO_CLK_c), .D(n5762));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4853_4854 (.Q(\REG.mem_50_5 ), .C(FIFO_CLK_c), .D(n5761));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4850_4851 (.Q(\REG.mem_50_4 ), .C(FIFO_CLK_c), .D(n5760));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4847_4848 (.Q(\REG.mem_50_3 ), .C(FIFO_CLK_c), .D(n5759));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4844_4845 (.Q(\REG.mem_50_2 ), .C(FIFO_CLK_c), .D(n5758));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4841_4842 (.Q(\REG.mem_50_1 ), .C(FIFO_CLK_c), .D(n5757));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY wr_addr_r_6__I_0_add_2_2 (.CI(VCC_net), .I0(wr_addr_r[0]), 
            .I1(rp_sync_w[0]), .CO(n10096));
    SB_LUT4 i9334_3_lut (.I0(\REG.mem_14_4 ), .I1(\REG.mem_15_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11172));
    defparam i9334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_8_lut (.I0(rd_sig_diff0_w[5]), .I1(wp_sync2_r[6]), 
            .I2(n1[6]), .I3(n10095), .O(n10873)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_7_lut (.I0(GND_net), .I1(wp_sync_w[5]), 
            .I2(n1[5]), .I3(n10094), .O(rd_sig_diff0_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9333_3_lut (.I0(\REG.mem_12_4 ), .I1(\REG.mem_13_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11171));
    defparam i9333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10011_3_lut (.I0(\REG.mem_0_14 ), .I1(\REG.mem_1_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11849));
    defparam i10011_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rd_addr_r_6__I_0_151_4 (.CI(n10140), .I0(rd_addr_r_c[2]), .I1(GND_net), 
            .CO(n10141));
    SB_DFF \REG.out_buffer__i14  (.Q(\fifo_data_out[14] ), .C(SLM_CLK_c), 
           .D(n10582));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i15  (.Q(\fifo_data_out[15] ), .C(SLM_CLK_c), 
           .D(n10588));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF i4838_4839 (.Q(\REG.mem_50_0 ), .C(FIFO_CLK_c), .D(n5753));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4787_4788 (.Q(\REG.mem_49_15 ), .C(FIFO_CLK_c), .D(n5752));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4784_4785 (.Q(\REG.mem_49_14 ), .C(FIFO_CLK_c), .D(n5751));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4781_4782 (.Q(\REG.mem_49_13 ), .C(FIFO_CLK_c), .D(n5750));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4778_4779 (.Q(\REG.mem_49_12 ), .C(FIFO_CLK_c), .D(n5749));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4775_4776 (.Q(\REG.mem_49_11 ), .C(FIFO_CLK_c), .D(n5748));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4772_4773 (.Q(\REG.mem_49_10 ), .C(FIFO_CLK_c), .D(n5747));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4769_4770 (.Q(\REG.mem_49_9 ), .C(FIFO_CLK_c), .D(n5746));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4766_4767 (.Q(\REG.mem_49_8 ), .C(FIFO_CLK_c), .D(n5745));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4763_4764 (.Q(\REG.mem_49_7 ), .C(FIFO_CLK_c), .D(n5744));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4760_4761 (.Q(\REG.mem_49_6 ), .C(FIFO_CLK_c), .D(n5743));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4757_4758 (.Q(\REG.mem_49_5 ), .C(FIFO_CLK_c), .D(n5742));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4754_4755 (.Q(\REG.mem_49_4 ), .C(FIFO_CLK_c), .D(n5741));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10012_3_lut (.I0(\REG.mem_2_14 ), .I1(\REG.mem_3_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11850));
    defparam i10012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_6__I_0_151_3_lut (.I0(GND_net), .I1(rd_addr_r_c[1]), 
            .I2(GND_net), .I3(n10139), .O(rd_addr_p1_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10015_3_lut (.I0(\REG.mem_6_14 ), .I1(\REG.mem_7_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11853));
    defparam i10015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10014_3_lut (.I0(\REG.mem_4_14 ), .I1(\REG.mem_5_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11852));
    defparam i10014_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rd_addr_r_6__I_0_151_3 (.CI(n10139), .I0(rd_addr_r_c[1]), .I1(GND_net), 
            .CO(n10140));
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_7 (.CI(n10094), .I0(wp_sync_w[5]), 
            .I1(n1[5]), .CO(n10095));
    SB_DFF i4751_4752 (.Q(\REG.mem_49_3 ), .C(FIFO_CLK_c), .D(n5740));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4748_4749 (.Q(\REG.mem_49_2 ), .C(FIFO_CLK_c), .D(n5739));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4745_4746 (.Q(\REG.mem_49_1 ), .C(FIFO_CLK_c), .D(n5738));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4742_4743 (.Q(\REG.mem_49_0 ), .C(FIFO_CLK_c), .D(n5737));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4691_4692 (.Q(\REG.mem_48_15 ), .C(FIFO_CLK_c), .D(n5736));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4688_4689 (.Q(\REG.mem_48_14 ), .C(FIFO_CLK_c), .D(n5735));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4685_4686 (.Q(\REG.mem_48_13 ), .C(FIFO_CLK_c), .D(n5734));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4682_4683 (.Q(\REG.mem_48_12 ), .C(FIFO_CLK_c), .D(n5733));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4679_4680 (.Q(\REG.mem_48_11 ), .C(FIFO_CLK_c), .D(n5732));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4676_4677 (.Q(\REG.mem_48_10 ), .C(FIFO_CLK_c), .D(n5731));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4673_4674 (.Q(\REG.mem_48_9 ), .C(FIFO_CLK_c), .D(n5730));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4670_4671 (.Q(\REG.mem_48_8 ), .C(FIFO_CLK_c), .D(n5729));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4667_4668 (.Q(\REG.mem_48_7 ), .C(FIFO_CLK_c), .D(n5728));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4664_4665 (.Q(\REG.mem_48_6 ), .C(FIFO_CLK_c), .D(n5727));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4661_4662 (.Q(\REG.mem_48_5 ), .C(FIFO_CLK_c), .D(n5726));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9171_3_lut (.I0(n12446), .I1(n12386), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11009));
    defparam i9171_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i4658_4659 (.Q(\REG.mem_48_4 ), .C(FIFO_CLK_c), .D(n5725));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4655_4656 (.Q(\REG.mem_48_3 ), .C(FIFO_CLK_c), .D(n5724));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_6_lut (.I0(rd_sig_diff0_w[3]), .I1(wp_sync_w[4]), 
            .I2(n1[4]), .I3(n10093), .O(n10877)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_6_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 n13133_bdd_4_lut (.I0(n13133), .I1(\REG.mem_9_15 ), .I2(\REG.mem_8_15 ), 
            .I3(rd_addr_r_c[1]), .O(n13136));
    defparam n13133_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11750 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_7 ), 
            .I2(\REG.mem_31_7 ), .I3(rd_addr_r_c[1]), .O(n13847));
    defparam rd_addr_r_0__bdd_4_lut_11750.LUT_INIT = 16'he4aa;
    SB_DFF i4652_4653 (.Q(\REG.mem_48_2 ), .C(FIFO_CLK_c), .D(n5723));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4649_4650 (.Q(\REG.mem_48_1 ), .C(FIFO_CLK_c), .D(n5722));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4646_4647 (.Q(\REG.mem_48_0 ), .C(FIFO_CLK_c), .D(n5721));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4595_4596 (.Q(\REG.mem_47_15 ), .C(FIFO_CLK_c), .D(n5720));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13847_bdd_4_lut (.I0(n13847), .I1(\REG.mem_29_7 ), .I2(\REG.mem_28_7 ), 
            .I3(rd_addr_r_c[1]), .O(n13850));
    defparam n13847_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4592_4593 (.Q(\REG.mem_47_14 ), .C(FIFO_CLK_c), .D(n5719));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i77_78 (.Q(\REG.mem_0_13 ), .C(FIFO_CLK_c), .D(n4926));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i80_81 (.Q(\REG.mem_0_14 ), .C(FIFO_CLK_c), .D(n4925));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9172_3_lut (.I0(n12368), .I1(n12350), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11010));
    defparam i9172_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i4589_4590 (.Q(\REG.mem_47_13 ), .C(FIFO_CLK_c), .D(n5718));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4586_4587 (.Q(\REG.mem_47_12 ), .C(FIFO_CLK_c), .D(n5717));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4583_4584 (.Q(\REG.mem_47_11 ), .C(FIFO_CLK_c), .D(n5716));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4580_4581 (.Q(\REG.mem_47_10 ), .C(FIFO_CLK_c), .D(n5715));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4577_4578 (.Q(\REG.mem_47_9 ), .C(FIFO_CLK_c), .D(n5714));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4574_4575 (.Q(\REG.mem_47_8 ), .C(FIFO_CLK_c), .D(n5713));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4571_4572 (.Q(\REG.mem_47_7 ), .C(FIFO_CLK_c), .D(n5712));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4568_4569 (.Q(\REG.mem_47_6 ), .C(FIFO_CLK_c), .D(n5711));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4565_4566 (.Q(\REG.mem_47_5 ), .C(FIFO_CLK_c), .D(n5710));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4562_4563 (.Q(\REG.mem_47_4 ), .C(FIFO_CLK_c), .D(n5709));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4559_4560 (.Q(\REG.mem_47_3 ), .C(FIFO_CLK_c), .D(n5708));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4556_4557 (.Q(\REG.mem_47_2 ), .C(FIFO_CLK_c), .D(n5707));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4553_4554 (.Q(\REG.mem_47_1 ), .C(FIFO_CLK_c), .D(n5706));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4550_4551 (.Q(\REG.mem_47_0 ), .C(FIFO_CLK_c), .D(n5705));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4499_4500 (.Q(\REG.mem_46_15 ), .C(FIFO_CLK_c), .D(n5704));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4496_4497 (.Q(\REG.mem_46_14 ), .C(FIFO_CLK_c), .D(n5703));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10627 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_0 ), 
            .I2(\REG.mem_63_0 ), .I3(rd_addr_r_c[1]), .O(n12479));
    defparam rd_addr_r_0__bdd_4_lut_10627.LUT_INIT = 16'he4aa;
    SB_DFF i83_84 (.Q(\REG.mem_0_15 ), .C(FIFO_CLK_c), .D(n4924));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12479_bdd_4_lut (.I0(n12479), .I1(\REG.mem_61_0 ), .I2(\REG.mem_60_0 ), 
            .I3(rd_addr_r_c[1]), .O(n12482));
    defparam n12479_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut (.I0(rd_addr_r_c[2]), .I1(n12422), .I2(n12380), 
            .I3(rd_addr_r_c[3]), .O(n13841));
    defparam rd_addr_r_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11150 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_12 ), 
            .I2(\REG.mem_31_12 ), .I3(rd_addr_r_c[1]), .O(n13127));
    defparam rd_addr_r_0__bdd_4_lut_11150.LUT_INIT = 16'he4aa;
    SB_DFF i4493_4494 (.Q(\REG.mem_46_13 ), .C(FIFO_CLK_c), .D(n5702));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9174_3_lut (.I0(n12338), .I1(n13814), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11012));
    defparam i9174_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i4490_4491 (.Q(\REG.mem_46_12 ), .C(FIFO_CLK_c), .D(n5701));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4487_4488 (.Q(\REG.mem_46_11 ), .C(FIFO_CLK_c), .D(n5700));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13841_bdd_4_lut (.I0(n13841), .I1(n12506), .I2(n12620), .I3(rd_addr_r_c[3]), 
            .O(n11401));
    defparam n13841_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4484_4485 (.Q(\REG.mem_46_10 ), .C(FIFO_CLK_c), .D(n5699));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3985_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_27_6 ), .O(n5368));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3985_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i4481_4482 (.Q(\REG.mem_46_9 ), .C(FIFO_CLK_c), .D(n5698));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13127_bdd_4_lut (.I0(n13127), .I1(\REG.mem_29_12 ), .I2(\REG.mem_28_12 ), 
            .I3(rd_addr_r_c[1]), .O(n13130));
    defparam n13127_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4478_4479 (.Q(\REG.mem_46_8 ), .C(FIFO_CLK_c), .D(n5697));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4475_4476 (.Q(\REG.mem_46_7 ), .C(FIFO_CLK_c), .D(n5696));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4472_4473 (.Q(\REG.mem_46_6 ), .C(FIFO_CLK_c), .D(n5695));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11145 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_3 ), 
            .I2(\REG.mem_55_3 ), .I3(rd_addr_r_c[1]), .O(n13121));
    defparam rd_addr_r_0__bdd_4_lut_11145.LUT_INIT = 16'he4aa;
    SB_DFF i4469_4470 (.Q(\REG.mem_46_5 ), .C(FIFO_CLK_c), .D(n5694));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4466_4467 (.Q(\REG.mem_46_4 ), .C(FIFO_CLK_c), .D(n5693));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4463_4464 (.Q(\REG.mem_46_3 ), .C(FIFO_CLK_c), .D(n5692));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4460_4461 (.Q(\REG.mem_46_2 ), .C(FIFO_CLK_c), .D(n5691));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4457_4458 (.Q(\REG.mem_46_1 ), .C(FIFO_CLK_c), .D(n5690));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4454_4455 (.Q(\REG.mem_46_0 ), .C(FIFO_CLK_c), .D(n5689));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4403_4404 (.Q(\REG.mem_45_15 ), .C(FIFO_CLK_c), .D(n5688));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4400_4401 (.Q(\REG.mem_45_14 ), .C(FIFO_CLK_c), .D(n5687));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4397_4398 (.Q(\REG.mem_45_13 ), .C(FIFO_CLK_c), .D(n5686));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4394_4395 (.Q(\REG.mem_45_12 ), .C(FIFO_CLK_c), .D(n5685));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4391_4392 (.Q(\REG.mem_45_11 ), .C(FIFO_CLK_c), .D(n5684));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4388_4389 (.Q(\REG.mem_45_10 ), .C(FIFO_CLK_c), .D(n5683));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4385_4386 (.Q(\REG.mem_45_9 ), .C(FIFO_CLK_c), .D(n5682));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4382_4383 (.Q(\REG.mem_45_8 ), .C(FIFO_CLK_c), .D(n5681));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4379_4380 (.Q(\REG.mem_45_7 ), .C(FIFO_CLK_c), .D(n5680));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4376_4377 (.Q(\REG.mem_45_6 ), .C(FIFO_CLK_c), .D(n5679));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut (.I0(rd_addr_r_c[1]), .I1(n11861), .I2(n11862), 
            .I3(rd_addr_r_c[2]), .O(n13835));
    defparam rd_addr_r_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n13121_bdd_4_lut (.I0(n13121), .I1(\REG.mem_53_3 ), .I2(\REG.mem_52_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11119));
    defparam n13121_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13835_bdd_4_lut (.I0(n13835), .I1(n11859), .I2(n11858), .I3(rd_addr_r_c[2]), 
            .O(n11025));
    defparam n13835_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4373_4374 (.Q(\REG.mem_45_5 ), .C(FIFO_CLK_c), .D(n5678));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11745 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_6 ), 
            .I2(\REG.mem_39_6 ), .I3(rd_addr_r_c[1]), .O(n13829));
    defparam rd_addr_r_0__bdd_4_lut_11745.LUT_INIT = 16'he4aa;
    SB_LUT4 i3984_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_27_5 ), .O(n5367));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3984_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3983_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_27_4 ), .O(n5366));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3983_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10742 (.I0(rd_addr_r_c[1]), .I1(n11897), 
            .I2(n11898), .I3(rd_addr_r_c[2]), .O(n12467));
    defparam rd_addr_r_1__bdd_4_lut_10742.LUT_INIT = 16'he4aa;
    SB_LUT4 n13829_bdd_4_lut (.I0(n13829), .I1(\REG.mem_37_6 ), .I2(\REG.mem_36_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11407));
    defparam n13829_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12467_bdd_4_lut (.I0(n12467), .I1(n11886), .I2(n11885), .I3(rd_addr_r_c[2]), 
            .O(n12470));
    defparam n12467_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4370_4371 (.Q(\REG.mem_45_4 ), .C(FIFO_CLK_c), .D(n5677));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11140 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_11 ), 
            .I2(\REG.mem_31_11 ), .I3(rd_addr_r_c[1]), .O(n13115));
    defparam rd_addr_r_0__bdd_4_lut_11140.LUT_INIT = 16'he4aa;
    SB_DFF i4367_4368 (.Q(\REG.mem_45_3 ), .C(FIFO_CLK_c), .D(n5676));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13115_bdd_4_lut (.I0(n13115), .I1(\REG.mem_29_11 ), .I2(\REG.mem_28_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11668));
    defparam n13115_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10607 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_5 ), 
            .I2(\REG.mem_43_5 ), .I3(rd_addr_r_c[1]), .O(n12461));
    defparam rd_addr_r_0__bdd_4_lut_10607.LUT_INIT = 16'he4aa;
    SB_DFF i4364_4365 (.Q(\REG.mem_45_2 ), .C(FIFO_CLK_c), .D(n5675));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4361_4362 (.Q(\REG.mem_45_1 ), .C(FIFO_CLK_c), .D(n5674));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4358_4359 (.Q(\REG.mem_45_0 ), .C(FIFO_CLK_c), .D(n5673));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wr_grey_sync_r__i6 (.Q(wr_grey_sync_r[6]), .C(FIFO_CLK_c), .D(n5672));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFF i4307_4308 (.Q(\REG.mem_44_15 ), .C(FIFO_CLK_c), .D(n5671));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4304_4305 (.Q(\REG.mem_44_14 ), .C(FIFO_CLK_c), .D(n5670));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4301_4302 (.Q(\REG.mem_44_13 ), .C(FIFO_CLK_c), .D(n5669));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4298_4299 (.Q(\REG.mem_44_12 ), .C(FIFO_CLK_c), .D(n5668));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4295_4296 (.Q(\REG.mem_44_11 ), .C(FIFO_CLK_c), .D(n5666));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4292_4293 (.Q(\REG.mem_44_10 ), .C(FIFO_CLK_c), .D(n5665));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4289_4290 (.Q(\REG.mem_44_9 ), .C(FIFO_CLK_c), .D(n5664));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4286_4287 (.Q(\REG.mem_44_8 ), .C(FIFO_CLK_c), .D(n5662));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4283_4284 (.Q(\REG.mem_44_7 ), .C(FIFO_CLK_c), .D(n5661));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_4__bdd_4_lut (.I0(rd_addr_r_c[4]), .I1(n11392), .I2(n11401), 
            .I3(rd_addr_r_c[5]), .O(n13823));
    defparam rd_addr_r_4__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11135 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_1 ), 
            .I2(\REG.mem_55_1 ), .I3(rd_addr_r_c[1]), .O(n13109));
    defparam rd_addr_r_0__bdd_4_lut_11135.LUT_INIT = 16'he4aa;
    SB_LUT4 i3982_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_27_3 ), .O(n5365));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3982_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13109_bdd_4_lut (.I0(n13109), .I1(\REG.mem_53_1 ), .I2(\REG.mem_52_1 ), 
            .I3(rd_addr_r_c[1]), .O(n13112));
    defparam n13109_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3981_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_27_2 ), .O(n5364));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3981_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3980_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_27_1 ), .O(n5363));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3980_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i4280_4281 (.Q(\REG.mem_44_6 ), .C(FIFO_CLK_c), .D(n5660));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4277_4278 (.Q(\REG.mem_44_5 ), .C(FIFO_CLK_c), .D(n5659));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4274_4275 (.Q(\REG.mem_44_4 ), .C(FIFO_CLK_c), .D(n5658));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4271_4272 (.Q(\REG.mem_44_3 ), .C(FIFO_CLK_c), .D(n5657));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4268_4269 (.Q(\REG.mem_44_2 ), .C(FIFO_CLK_c), .D(n5656));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4265_4266 (.Q(\REG.mem_44_1 ), .C(FIFO_CLK_c), .D(n5655));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4262_4263 (.Q(\REG.mem_44_0 ), .C(FIFO_CLK_c), .D(n5654));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4211_4212 (.Q(\REG.mem_43_15 ), .C(FIFO_CLK_c), .D(n5653));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4208_4209 (.Q(\REG.mem_43_14 ), .C(FIFO_CLK_c), .D(n5652));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4205_4206 (.Q(\REG.mem_43_13 ), .C(FIFO_CLK_c), .D(n5651));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4202_4203 (.Q(\REG.mem_43_12 ), .C(FIFO_CLK_c), .D(n5650));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4199_4200 (.Q(\REG.mem_43_11 ), .C(FIFO_CLK_c), .D(n5649));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4196_4197 (.Q(\REG.mem_43_10 ), .C(FIFO_CLK_c), .D(n5648));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4193_4194 (.Q(\REG.mem_43_9 ), .C(FIFO_CLK_c), .D(n5647));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4190_4191 (.Q(\REG.mem_43_8 ), .C(FIFO_CLK_c), .D(n5646));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4187_4188 (.Q(\REG.mem_43_7 ), .C(FIFO_CLK_c), .D(n5645));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4184_4185 (.Q(\REG.mem_43_6 ), .C(FIFO_CLK_c), .D(n5644));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3979_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_27_0 ), .O(n5362));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3979_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12461_bdd_4_lut (.I0(n12461), .I1(\REG.mem_41_5 ), .I2(\REG.mem_40_5 ), 
            .I3(rd_addr_r_c[1]), .O(n12464));
    defparam n12461_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13823_bdd_4_lut (.I0(n13823), .I1(n11383), .I2(n12320), .I3(rd_addr_r_c[5]), 
            .O(\REG.out_raw_31__N_559 [9]));
    defparam n13823_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_6 (.CI(n10093), .I0(wp_sync_w[4]), 
            .I1(n1[4]), .CO(n10094));
    SB_LUT4 i4010_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_28_15 ), .O(n5393));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4010_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4009_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_28_14 ), .O(n5392));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4009_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4008_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_28_13 ), .O(n5391));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4008_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_5_lut (.I0(GND_net), .I1(wp_sync_w[3]), 
            .I2(n1[3]), .I3(n10092), .O(rd_sig_diff0_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11730 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_1 ), 
            .I2(\REG.mem_23_1 ), .I3(rd_addr_r_c[1]), .O(n13817));
    defparam rd_addr_r_0__bdd_4_lut_11730.LUT_INIT = 16'he4aa;
    SB_LUT4 i4007_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_28_12 ), .O(n5390));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4007_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_6__I_0_151_2_lut (.I0(GND_net), .I1(rd_addr_r[0]), 
            .I2(GND_net), .I3(VCC_net), .O(\rd_addr_p1_w[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_5 (.CI(n10092), .I0(wp_sync_w[3]), 
            .I1(n1[3]), .CO(n10093));
    SB_LUT4 n13817_bdd_4_lut (.I0(n13817), .I1(\REG.mem_21_1 ), .I2(\REG.mem_20_1 ), 
            .I3(rd_addr_r_c[1]), .O(n11419));
    defparam n13817_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11130 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_11 ), 
            .I2(\REG.mem_35_11 ), .I3(rd_addr_r_c[1]), .O(n13103));
    defparam rd_addr_r_0__bdd_4_lut_11130.LUT_INIT = 16'he4aa;
    SB_DFF i4181_4182 (.Q(\REG.mem_43_5 ), .C(FIFO_CLK_c), .D(n5643));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13103_bdd_4_lut (.I0(n13103), .I1(\REG.mem_33_11 ), .I2(\REG.mem_32_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11674));
    defparam n13103_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4178_4179 (.Q(\REG.mem_43_4 ), .C(FIFO_CLK_c), .D(n5642));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4175_4176 (.Q(\REG.mem_43_3 ), .C(FIFO_CLK_c), .D(n5641));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4172_4173 (.Q(\REG.mem_43_2 ), .C(FIFO_CLK_c), .D(n5640));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4169_4170 (.Q(\REG.mem_43_1 ), .C(FIFO_CLK_c), .D(n5639));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4166_4167 (.Q(\REG.mem_43_0 ), .C(FIFO_CLK_c), .D(n5638));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4115_4116 (.Q(\REG.mem_42_15 ), .C(FIFO_CLK_c), .D(n5637));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4112_4113 (.Q(\REG.mem_42_14 ), .C(FIFO_CLK_c), .D(n5636));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4109_4110 (.Q(\REG.mem_42_13 ), .C(FIFO_CLK_c), .D(n5635));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4106_4107 (.Q(\REG.mem_42_12 ), .C(FIFO_CLK_c), .D(n5634));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4103_4104 (.Q(\REG.mem_42_11 ), .C(FIFO_CLK_c), .D(n5633));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4100_4101 (.Q(\REG.mem_42_10 ), .C(FIFO_CLK_c), .D(n5632));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4097_4098 (.Q(\REG.mem_42_9 ), .C(FIFO_CLK_c), .D(n5631));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4094_4095 (.Q(\REG.mem_42_8 ), .C(FIFO_CLK_c), .D(n5630));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4091_4092 (.Q(\REG.mem_42_7 ), .C(FIFO_CLK_c), .D(n5629));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF \genblk16.rd_prev_r_132  (.Q(\genblk16.rd_prev_r ), .C(SLM_CLK_c), 
           .D(n4916));   // src/fifo_dc_32_lut_gen.v(751[29] 761[32])
    SB_LUT4 i4006_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_28_11 ), .O(n5389));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4006_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10539 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_15 ), 
            .I2(\REG.mem_43_15 ), .I3(rd_addr_r_c[1]), .O(n12389));
    defparam rd_addr_r_0__bdd_4_lut_10539.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10642 (.I0(rd_addr_r_c[2]), .I1(n11302), 
            .I2(n12434), .I3(rd_addr_r_c[3]), .O(n12455));
    defparam rd_addr_r_2__bdd_4_lut_10642.LUT_INIT = 16'he4aa;
    SB_LUT4 n12455_bdd_4_lut (.I0(n12455), .I1(n11230), .I2(n12416), .I3(rd_addr_r_c[3]), 
            .O(n12458));
    defparam n12455_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10592 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_6 ), 
            .I2(\REG.mem_31_6 ), .I3(rd_addr_r_c[1]), .O(n12449));
    defparam rd_addr_r_0__bdd_4_lut_10592.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11720 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_2 ), 
            .I2(\REG.mem_23_2 ), .I3(rd_addr_r_c[1]), .O(n13811));
    defparam rd_addr_r_0__bdd_4_lut_11720.LUT_INIT = 16'he4aa;
    SB_LUT4 n12449_bdd_4_lut (.I0(n12449), .I1(\REG.mem_29_6 ), .I2(\REG.mem_28_6 ), 
            .I3(rd_addr_r_c[1]), .O(n12452));
    defparam n12449_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11125 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_11 ), 
            .I2(\REG.mem_39_11 ), .I3(rd_addr_r_c[1]), .O(n13097));
    defparam rd_addr_r_0__bdd_4_lut_11125.LUT_INIT = 16'he4aa;
    SB_LUT4 n13097_bdd_4_lut (.I0(n13097), .I1(\REG.mem_37_11 ), .I2(\REG.mem_36_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11677));
    defparam n13097_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i167_168 (.Q(\REG.mem_1_11 ), .C(FIFO_CLK_c), .D(n4915));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i152_153 (.Q(\REG.mem_1_6 ), .C(FIFO_CLK_c), .D(n4914));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4088_4089 (.Q(\REG.mem_42_6 ), .C(FIFO_CLK_c), .D(n5628));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4085_4086 (.Q(\REG.mem_42_5 ), .C(FIFO_CLK_c), .D(n5627));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4082_4083 (.Q(\REG.mem_42_4 ), .C(FIFO_CLK_c), .D(n5626));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4079_4080 (.Q(\REG.mem_42_3 ), .C(FIFO_CLK_c), .D(n5625));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4076_4077 (.Q(\REG.mem_42_2 ), .C(FIFO_CLK_c), .D(n5624));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4073_4074 (.Q(\REG.mem_42_1 ), .C(FIFO_CLK_c), .D(n5623));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4070_4071 (.Q(\REG.mem_42_0 ), .C(FIFO_CLK_c), .D(n5622));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4019_4020 (.Q(\REG.mem_41_15 ), .C(FIFO_CLK_c), .D(n5621));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4016_4017 (.Q(\REG.mem_41_14 ), .C(FIFO_CLK_c), .D(n5620));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4013_4014 (.Q(\REG.mem_41_13 ), .C(FIFO_CLK_c), .D(n5619));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4010_4011 (.Q(\REG.mem_41_12 ), .C(FIFO_CLK_c), .D(n5618));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4007_4008 (.Q(\REG.mem_41_11 ), .C(FIFO_CLK_c), .D(n5617));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4004_4005 (.Q(\REG.mem_41_10 ), .C(FIFO_CLK_c), .D(n5616));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4001_4002 (.Q(\REG.mem_41_9 ), .C(FIFO_CLK_c), .D(n5615));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3998_3999 (.Q(\REG.mem_41_8 ), .C(FIFO_CLK_c), .D(n5614));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3995_3996 (.Q(\REG.mem_41_7 ), .C(FIFO_CLK_c), .D(n5613));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4005_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_28_10 ), .O(n5388));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4005_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4004_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_28_9 ), .O(n5387));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4004_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13811_bdd_4_lut (.I0(n13811), .I1(\REG.mem_21_2 ), .I2(\REG.mem_20_2 ), 
            .I3(rd_addr_r_c[1]), .O(n13814));
    defparam n13811_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11510 (.I0(rd_addr_r_c[2]), .I1(n12830), 
            .I2(n12770), .I3(rd_addr_r_c[3]), .O(n13091));
    defparam rd_addr_r_2__bdd_4_lut_11510.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10582 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_2 ), 
            .I2(\REG.mem_3_2 ), .I3(rd_addr_r_c[1]), .O(n12443));
    defparam rd_addr_r_0__bdd_4_lut_10582.LUT_INIT = 16'he4aa;
    SB_LUT4 n12443_bdd_4_lut (.I0(n12443), .I1(\REG.mem_1_2 ), .I2(\REG.mem_0_2 ), 
            .I3(rd_addr_r_c[1]), .O(n12446));
    defparam n12443_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i170_171 (.Q(\REG.mem_1_12 ), .C(FIFO_CLK_c), .D(n4912));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3992_3993 (.Q(\REG.mem_41_6 ), .C(FIFO_CLK_c), .D(n5612));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3989_3990 (.Q(\REG.mem_41_5 ), .C(FIFO_CLK_c), .D(n5611));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3986_3987 (.Q(\REG.mem_41_4 ), .C(FIFO_CLK_c), .D(n5610));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3983_3984 (.Q(\REG.mem_41_3 ), .C(FIFO_CLK_c), .D(n5609));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3980_3981 (.Q(\REG.mem_41_2 ), .C(FIFO_CLK_c), .D(n5608));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3977_3978 (.Q(\REG.mem_41_1 ), .C(FIFO_CLK_c), .D(n5607));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3974_3975 (.Q(\REG.mem_41_0 ), .C(FIFO_CLK_c), .D(n5606));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3923_3924 (.Q(\REG.mem_40_15 ), .C(FIFO_CLK_c), .D(n5605));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3920_3921 (.Q(\REG.mem_40_14 ), .C(FIFO_CLK_c), .D(n5604));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3917_3918 (.Q(\REG.mem_40_13 ), .C(FIFO_CLK_c), .D(n5603));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3914_3915 (.Q(\REG.mem_40_12 ), .C(FIFO_CLK_c), .D(n5602));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3911_3912 (.Q(\REG.mem_40_11 ), .C(FIFO_CLK_c), .D(n5601));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3908_3909 (.Q(\REG.mem_40_10 ), .C(FIFO_CLK_c), .D(n5600));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3905_3906 (.Q(\REG.mem_40_9 ), .C(FIFO_CLK_c), .D(n5599));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3902_3903 (.Q(\REG.mem_40_8 ), .C(FIFO_CLK_c), .D(n5598));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3899_3900 (.Q(\REG.mem_40_7 ), .C(FIFO_CLK_c), .D(n5597));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9393_3_lut (.I0(\REG.mem_24_9 ), .I1(\REG.mem_25_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11231));
    defparam i9393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13091_bdd_4_lut (.I0(n13091), .I1(n12854), .I2(n12914), .I3(rd_addr_r_c[3]), 
            .O(n13094));
    defparam n13091_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11715 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_14 ), 
            .I2(\REG.mem_63_14 ), .I3(rd_addr_r_c[1]), .O(n13805));
    defparam rd_addr_r_0__bdd_4_lut_11715.LUT_INIT = 16'he4aa;
    SB_LUT4 i4003_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_28_8 ), .O(n5386));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4003_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY rd_addr_r_6__I_0_151_2 (.CI(VCC_net), .I0(rd_addr_r[0]), .I1(GND_net), 
            .CO(n10139));
    SB_DFF i155_156 (.Q(\REG.mem_1_7 ), .C(FIFO_CLK_c), .D(n4905));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9394_3_lut (.I0(\REG.mem_26_9 ), .I1(\REG.mem_27_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11232));
    defparam i9394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13805_bdd_4_lut (.I0(n13805), .I1(\REG.mem_61_14 ), .I2(\REG.mem_60_14 ), 
            .I3(rd_addr_r_c[1]), .O(n10996));
    defparam n13805_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF wp_sync2_r__i0 (.Q(wp_sync2_r[0]), .C(SLM_CLK_c), .D(n4904));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_LUT4 i4002_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_28_7 ), .O(n5385));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4002_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF wp_sync1_r__i0 (.Q(wp_sync1_r[0]), .C(SLM_CLK_c), .D(n4903));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF i173_174 (.Q(\REG.mem_1_13 ), .C(FIFO_CLK_c), .D(n4902));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rd_addr_r__i0 (.Q(rd_addr_r[0]), .C(SLM_CLK_c), .D(n4901));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF i158_159 (.Q(\REG.mem_1_8 ), .C(FIFO_CLK_c), .D(n4900));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync2_r__i0 (.Q(rp_sync2_r[0]), .C(FIFO_CLK_c), .D(n4899));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF i3896_3897 (.Q(\REG.mem_40_6 ), .C(FIFO_CLK_c), .D(n5596));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11170 (.I0(rd_addr_r_c[3]), .I1(n11567), 
            .I2(n11568), .I3(rd_addr_r_c[4]), .O(n13085));
    defparam rd_addr_r_3__bdd_4_lut_11170.LUT_INIT = 16'he4aa;
    SB_DFF i3893_3894 (.Q(\REG.mem_40_5 ), .C(FIFO_CLK_c), .D(n5595));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3890_3891 (.Q(\REG.mem_40_4 ), .C(FIFO_CLK_c), .D(n5594));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3887_3888 (.Q(\REG.mem_40_3 ), .C(FIFO_CLK_c), .D(n5593));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3884_3885 (.Q(\REG.mem_40_2 ), .C(FIFO_CLK_c), .D(n5592));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3881_3882 (.Q(\REG.mem_40_1 ), .C(FIFO_CLK_c), .D(n5591));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3878_3879 (.Q(\REG.mem_40_0 ), .C(FIFO_CLK_c), .D(n5590));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3827_3828 (.Q(\REG.mem_39_15 ), .C(FIFO_CLK_c), .D(n5589));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3824_3825 (.Q(\REG.mem_39_14 ), .C(FIFO_CLK_c), .D(n5588));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3821_3822 (.Q(\REG.mem_39_13 ), .C(FIFO_CLK_c), .D(n5587));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3818_3819 (.Q(\REG.mem_39_12 ), .C(FIFO_CLK_c), .D(n5586));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3815_3816 (.Q(\REG.mem_39_11 ), .C(FIFO_CLK_c), .D(n5585));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3812_3813 (.Q(\REG.mem_39_10 ), .C(FIFO_CLK_c), .D(n5584));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3809_3810 (.Q(\REG.mem_39_9 ), .C(FIFO_CLK_c), .D(n5583));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3806_3807 (.Q(\REG.mem_39_8 ), .C(FIFO_CLK_c), .D(n5582));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3803_3804 (.Q(\REG.mem_39_7 ), .C(FIFO_CLK_c), .D(n5581));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync1_r__i0 (.Q(rp_sync1_r[0]), .C(FIFO_CLK_c), .D(n4898));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_LUT4 rd_addr_r_3__bdd_4_lut (.I0(rd_addr_r_c[3]), .I1(n12680), .I2(n11022), 
            .I3(rd_addr_r_c[4]), .O(n13799));
    defparam rd_addr_r_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n13799_bdd_4_lut (.I0(n13799), .I1(n11019), .I2(n12674), .I3(rd_addr_r_c[4]), 
            .O(n13802));
    defparam n13799_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut (.I0(wr_sig_diff0_w[0]), .I1(wr_sig_diff0_w[1]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_23));   // src/fifo_dc_32_lut_gen.v(403[38:87])
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10577 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_1 ), 
            .I2(\REG.mem_15_1 ), .I3(rd_addr_r_c[1]), .O(n12431));
    defparam rd_addr_r_0__bdd_4_lut_10577.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut (.I0(DEBUG_5_c), .I1(wr_sig_diff0_w[3]), .I2(n6_adj_23), 
            .I3(wr_sig_diff0_w[2]), .O(n2_adj_22));   // src/fifo_dc_32_lut_gen.v(403[38:87])
    defparam i1_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 n12431_bdd_4_lut (.I0(n12431), .I1(\REG.mem_13_1 ), .I2(\REG.mem_12_1 ), 
            .I3(rd_addr_r_c[1]), .O(n12434));
    defparam n12431_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13085_bdd_4_lut (.I0(n13085), .I1(n11553), .I2(n13040), .I3(rd_addr_r_c[4]), 
            .O(n13088));
    defparam n13085_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11710 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_3 ), 
            .I2(\REG.mem_3_3 ), .I3(rd_addr_r_c[1]), .O(n13793));
    defparam rd_addr_r_0__bdd_4_lut_11710.LUT_INIT = 16'he4aa;
    SB_LUT4 n13793_bdd_4_lut (.I0(n13793), .I1(\REG.mem_1_3 ), .I2(\REG.mem_0_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11035));
    defparam n13793_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut (.I0(wr_sig_diff0_w[2]), .I1(wr_sig_diff0_w[1]), .I2(wr_sig_diff0_w[0]), 
            .I3(GND_net), .O(n10254));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9114_4_lut (.I0(dc32_fifo_almost_full), .I1(n10925), .I2(n10254), 
            .I3(wr_sig_diff0_w[3]), .O(n10951));
    defparam i9114_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11110 (.I0(rd_addr_r_c[3]), .I1(n13046), 
            .I2(n11559), .I3(rd_addr_r_c[4]), .O(n13079));
    defparam rd_addr_r_3__bdd_4_lut_11110.LUT_INIT = 16'he4aa;
    SB_LUT4 n13079_bdd_4_lut (.I0(n13079), .I1(n11550), .I2(n13034), .I3(rd_addr_r_c[4]), 
            .O(n13082));
    defparam n13079_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4001_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_28_6 ), .O(n5384));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4001_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3800_3801 (.Q(\REG.mem_39_6 ), .C(FIFO_CLK_c), .D(n5580));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3797_3798 (.Q(\REG.mem_39_5 ), .C(FIFO_CLK_c), .D(n5579));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4000_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_28_5 ), .O(n5383));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4000_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3794_3795 (.Q(\REG.mem_39_4 ), .C(FIFO_CLK_c), .D(n5578));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3791_3792 (.Q(\REG.mem_39_3 ), .C(FIFO_CLK_c), .D(n5577));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3788_3789 (.Q(\REG.mem_39_2 ), .C(FIFO_CLK_c), .D(n5576));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3785_3786 (.Q(\REG.mem_39_1 ), .C(FIFO_CLK_c), .D(n5575));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3782_3783 (.Q(\REG.mem_39_0 ), .C(FIFO_CLK_c), .D(n5573));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3731_3732 (.Q(\REG.mem_38_15 ), .C(FIFO_CLK_c), .D(n5572));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3728_3729 (.Q(\REG.mem_38_14 ), .C(FIFO_CLK_c), .D(n5571));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3725_3726 (.Q(\REG.mem_38_13 ), .C(FIFO_CLK_c), .D(n5570));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3722_3723 (.Q(\REG.mem_38_12 ), .C(FIFO_CLK_c), .D(n5569));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3719_3720 (.Q(\REG.mem_38_11 ), .C(FIFO_CLK_c), .D(n5568));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3716_3717 (.Q(\REG.mem_38_10 ), .C(FIFO_CLK_c), .D(n5567));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3713_3714 (.Q(\REG.mem_38_9 ), .C(FIFO_CLK_c), .D(n5566));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3710_3711 (.Q(\REG.mem_38_8 ), .C(FIFO_CLK_c), .D(n5565));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3707_3708 (.Q(\REG.mem_38_7 ), .C(FIFO_CLK_c), .D(n5564));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3999_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_28_4 ), .O(n5382));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3999_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3998_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_28_3 ), .O(n5381));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3998_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3997_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_28_2 ), .O(n5380));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3997_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3996_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_28_1 ), .O(n5379));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3996_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3995_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_28_0 ), .O(n5378));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3995_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4026_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_29_15 ), .O(n5409));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4026_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4025_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_29_14 ), .O(n5408));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4025_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12389_bdd_4_lut (.I0(n12389), .I1(\REG.mem_41_15 ), .I2(\REG.mem_40_15 ), 
            .I3(rd_addr_r_c[1]), .O(n12392));
    defparam n12389_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4024_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_29_13 ), .O(n5407));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4024_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4023_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_29_12 ), .O(n5406));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4023_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4022_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_29_11 ), .O(n5405));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4022_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4021_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_29_10 ), .O(n5404));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4021_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10499 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_5 ), 
            .I2(\REG.mem_47_5 ), .I3(rd_addr_r_c[1]), .O(n12341));
    defparam rd_addr_r_0__bdd_4_lut_10499.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11700 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_13 ), 
            .I2(\REG.mem_43_13 ), .I3(rd_addr_r_c[1]), .O(n13787));
    defparam rd_addr_r_0__bdd_4_lut_11700.LUT_INIT = 16'he4aa;
    SB_LUT4 n13787_bdd_4_lut (.I0(n13787), .I1(\REG.mem_41_13 ), .I2(\REG.mem_40_13 ), 
            .I3(rd_addr_r_c[1]), .O(n11440));
    defparam n13787_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4020_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_29_9 ), .O(n5403));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4020_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3704_3705 (.Q(\REG.mem_38_6 ), .C(FIFO_CLK_c), .D(n5563));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3701_3702 (.Q(\REG.mem_38_5 ), .C(FIFO_CLK_c), .D(n5562));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3698_3699 (.Q(\REG.mem_38_4 ), .C(FIFO_CLK_c), .D(n5561));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3695_3696 (.Q(\REG.mem_38_3 ), .C(FIFO_CLK_c), .D(n5560));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3692_3693 (.Q(\REG.mem_38_2 ), .C(FIFO_CLK_c), .D(n5559));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3689_3690 (.Q(\REG.mem_38_1 ), .C(FIFO_CLK_c), .D(n5558));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3686_3687 (.Q(\REG.mem_38_0 ), .C(FIFO_CLK_c), .D(n5556));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3635_3636 (.Q(\REG.mem_37_15 ), .C(FIFO_CLK_c), .D(n5555));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3632_3633 (.Q(\REG.mem_37_14 ), .C(FIFO_CLK_c), .D(n5554));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3629_3630 (.Q(\REG.mem_37_13 ), .C(FIFO_CLK_c), .D(n5553));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3626_3627 (.Q(\REG.mem_37_12 ), .C(FIFO_CLK_c), .D(n5552));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3623_3624 (.Q(\REG.mem_37_11 ), .C(FIFO_CLK_c), .D(n5551));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3620_3621 (.Q(\REG.mem_37_10 ), .C(FIFO_CLK_c), .D(n5550));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3617_3618 (.Q(\REG.mem_37_9 ), .C(FIFO_CLK_c), .D(n5549));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11155 (.I0(rd_addr_r_c[1]), .I1(n11504), 
            .I2(n11505), .I3(rd_addr_r_c[2]), .O(n13073));
    defparam rd_addr_r_1__bdd_4_lut_11155.LUT_INIT = 16'he4aa;
    SB_LUT4 n13073_bdd_4_lut (.I0(n13073), .I1(n11475), .I2(n11474), .I3(rd_addr_r_c[2]), 
            .O(n13076));
    defparam n13073_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11695 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_13 ), 
            .I2(\REG.mem_27_13 ), .I3(rd_addr_r_c[1]), .O(n13781));
    defparam rd_addr_r_0__bdd_4_lut_11695.LUT_INIT = 16'he4aa;
    SB_LUT4 i4019_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_29_8 ), .O(n5402));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4019_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13781_bdd_4_lut (.I0(n13781), .I1(\REG.mem_25_13 ), .I2(\REG.mem_24_13 ), 
            .I3(rd_addr_r_c[1]), .O(n13784));
    defparam n13781_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4018_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_29_7 ), .O(n5401));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4018_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \REG.out_raw__i16  (.Q(\REG.out_raw[15] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [15]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i15  (.Q(\REG.out_raw[14] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [14]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i14  (.Q(\REG.out_raw[13] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [13]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i13  (.Q(\REG.out_raw[12] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [12]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i12  (.Q(\REG.out_raw[11] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [11]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFF i3614_3615 (.Q(\REG.mem_37_8 ), .C(FIFO_CLK_c), .D(n5548));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3611_3612 (.Q(\REG.mem_37_7 ), .C(FIFO_CLK_c), .D(n5547));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3608_3609 (.Q(\REG.mem_37_6 ), .C(FIFO_CLK_c), .D(n5546));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3605_3606 (.Q(\REG.mem_37_5 ), .C(FIFO_CLK_c), .D(n5545));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3602_3603 (.Q(\REG.mem_37_4 ), .C(FIFO_CLK_c), .D(n5544));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3599_3600 (.Q(\REG.mem_37_3 ), .C(FIFO_CLK_c), .D(n5543));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3596_3597 (.Q(\REG.mem_37_2 ), .C(FIFO_CLK_c), .D(n5542));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3593_3594 (.Q(\REG.mem_37_1 ), .C(FIFO_CLK_c), .D(n5541));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3590_3591 (.Q(\REG.mem_37_0 ), .C(FIFO_CLK_c), .D(n5540));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11100 (.I0(rd_addr_r_c[1]), .I1(n11519), 
            .I2(n11520), .I3(rd_addr_r_c[2]), .O(n13067));
    defparam rd_addr_r_1__bdd_4_lut_11100.LUT_INIT = 16'he4aa;
    SB_LUT4 i4017_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_29_6 ), .O(n5400));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4017_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \REG.out_raw__i11  (.Q(\REG.out_raw[10] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [10]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i10  (.Q(\REG.out_raw[9] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [9]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i9  (.Q(\REG.out_raw[8] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [8]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFSR wr_grey_sync_r__i5 (.Q(wr_grey_sync_r[5]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[5]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFE \REG.out_raw__i8  (.Q(\REG.out_raw[7] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [7]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFSR wr_grey_sync_r__i4 (.Q(wr_grey_sync_r[4]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[4]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFE \REG.out_raw__i7  (.Q(\REG.out_raw[6] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [6]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFSR wr_grey_sync_r__i3 (.Q(wr_grey_sync_r[3]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[3]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFE \REG.out_raw__i6  (.Q(\REG.out_raw[5] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [5]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFSR wr_grey_sync_r__i2 (.Q(wr_grey_sync_r[2]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[2]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFE \REG.out_raw__i5  (.Q(\REG.out_raw[4] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [4]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFSR wr_grey_sync_r__i1 (.Q(wr_grey_sync_r[1]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[1]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFE \REG.out_raw__i4  (.Q(\REG.out_raw[3] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [3]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i3  (.Q(\REG.out_raw[2] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [2]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i2  (.Q(\REG.out_raw[1] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [1]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11690 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_2 ), 
            .I2(\REG.mem_43_2 ), .I3(rd_addr_r_c[1]), .O(n13775));
    defparam rd_addr_r_0__bdd_4_lut_11690.LUT_INIT = 16'he4aa;
    SB_LUT4 i4016_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_29_5 ), .O(n5399));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4016_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3539_3540 (.Q(\REG.mem_36_15 ), .C(FIFO_CLK_c), .D(n5526));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3536_3537 (.Q(\REG.mem_36_14 ), .C(FIFO_CLK_c), .D(n5525));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3533_3534 (.Q(\REG.mem_36_13 ), .C(FIFO_CLK_c), .D(n5524));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3530_3531 (.Q(\REG.mem_36_12 ), .C(FIFO_CLK_c), .D(n5523));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3527_3528 (.Q(\REG.mem_36_11 ), .C(FIFO_CLK_c), .D(n5522));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3524_3525 (.Q(\REG.mem_36_10 ), .C(FIFO_CLK_c), .D(n5521));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3521_3522 (.Q(\REG.mem_36_9 ), .C(FIFO_CLK_c), .D(n5520));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3518_3519 (.Q(\REG.mem_36_8 ), .C(FIFO_CLK_c), .D(n5519));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3515_3516 (.Q(\REG.mem_36_7 ), .C(FIFO_CLK_c), .D(n5518));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3512_3513 (.Q(\REG.mem_36_6 ), .C(FIFO_CLK_c), .D(n5517));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3509_3510 (.Q(\REG.mem_36_5 ), .C(FIFO_CLK_c), .D(n5516));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4015_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_29_4 ), .O(n5398));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4015_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10017_3_lut (.I0(\REG.mem_48_8 ), .I1(\REG.mem_49_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11855));
    defparam i10017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_141_8_lut (.I0(GND_net), .I1(wr_grey_sync_r[6]), 
            .I2(GND_net), .I3(n10138), .O(wr_addr_p1_w[6])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_4_lut (.I0(GND_net), .I1(wp_sync_w[2]), 
            .I2(n1[2]), .I3(n10091), .O(\rd_sig_diff0_w[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4014_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_29_3 ), .O(n5397));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4014_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3506_3507 (.Q(\REG.mem_36_4 ), .C(FIFO_CLK_c), .D(n5515));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3503_3504 (.Q(\REG.mem_36_3 ), .C(FIFO_CLK_c), .D(n5514));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3500_3501 (.Q(\REG.mem_36_2 ), .C(FIFO_CLK_c), .D(n5513));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3497_3498 (.Q(\REG.mem_36_1 ), .C(FIFO_CLK_c), .D(n5512));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3494_3495 (.Q(\REG.mem_36_0 ), .C(FIFO_CLK_c), .D(n5511));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3443_3444 (.Q(\REG.mem_35_15 ), .C(FIFO_CLK_c), .D(n5507));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4013_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_29_2 ), .O(n5396));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4013_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3440_3441 (.Q(\REG.mem_35_14 ), .C(FIFO_CLK_c), .D(n5506));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3437_3438 (.Q(\REG.mem_35_13 ), .C(FIFO_CLK_c), .D(n5505));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3434_3435 (.Q(\REG.mem_35_12 ), .C(FIFO_CLK_c), .D(n5504));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3431_3432 (.Q(\REG.mem_35_11 ), .C(FIFO_CLK_c), .D(n5503));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3428_3429 (.Q(\REG.mem_35_10 ), .C(FIFO_CLK_c), .D(n5502));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3425_3426 (.Q(\REG.mem_35_9 ), .C(FIFO_CLK_c), .D(n5501));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3422_3423 (.Q(\REG.mem_35_8 ), .C(FIFO_CLK_c), .D(n5500));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10018_3_lut (.I0(\REG.mem_50_8 ), .I1(\REG.mem_51_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11856));
    defparam i10018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13775_bdd_4_lut (.I0(n13775), .I1(\REG.mem_41_2 ), .I2(\REG.mem_40_2 ), 
            .I3(rd_addr_r_c[1]), .O(n13778));
    defparam n13775_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_4 (.CI(n10091), .I0(wp_sync_w[2]), 
            .I1(n1[2]), .CO(n10092));
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_3_lut (.I0(GND_net), .I1(wp_sync_w[1]), 
            .I2(n1[1]), .I3(n10090), .O(\rd_sig_diff0_w[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10027_3_lut (.I0(\REG.mem_54_8 ), .I1(\REG.mem_55_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11865));
    defparam i10027_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i3419_3420 (.Q(\REG.mem_35_7 ), .C(FIFO_CLK_c), .D(n5499));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3416_3417 (.Q(\REG.mem_35_6 ), .C(FIFO_CLK_c), .D(n5498));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3413_3414 (.Q(\REG.mem_35_5 ), .C(FIFO_CLK_c), .D(n5497));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3410_3411 (.Q(\REG.mem_35_4 ), .C(FIFO_CLK_c), .D(n5496));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3407_3408 (.Q(\REG.mem_35_3 ), .C(FIFO_CLK_c), .D(n5495));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3404_3405 (.Q(\REG.mem_35_2 ), .C(FIFO_CLK_c), .D(n5494));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3401_3402 (.Q(\REG.mem_35_1 ), .C(FIFO_CLK_c), .D(n5493));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3398_3399 (.Q(\REG.mem_35_0 ), .C(FIFO_CLK_c), .D(n5492));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3347_3348 (.Q(\REG.mem_34_15 ), .C(FIFO_CLK_c), .D(n5490));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3344_3345 (.Q(\REG.mem_34_14 ), .C(FIFO_CLK_c), .D(n5489));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3341_3342 (.Q(\REG.mem_34_13 ), .C(FIFO_CLK_c), .D(n5488));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3338_3339 (.Q(\REG.mem_34_12 ), .C(FIFO_CLK_c), .D(n5487));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3335_3336 (.Q(\REG.mem_34_11 ), .C(FIFO_CLK_c), .D(n5486));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3332_3333 (.Q(\REG.mem_34_10 ), .C(FIFO_CLK_c), .D(n5485));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3329_3330 (.Q(\REG.mem_34_9 ), .C(FIFO_CLK_c), .D(n5484));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4012_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_29_1 ), .O(n5395));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4012_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4011_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_29_0 ), .O(n5394));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4011_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4042_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_30_15 ), .O(n5425));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4042_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10026_3_lut (.I0(\REG.mem_52_8 ), .I1(\REG.mem_53_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11864));
    defparam i10026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4041_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_30_14 ), .O(n5424));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4041_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4040_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_30_13 ), .O(n5423));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4040_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4039_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_30_12 ), .O(n5422));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4039_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4038_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_30_11 ), .O(n5421));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4038_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11735 (.I0(rd_addr_r_c[1]), .I1(n11441), 
            .I2(n11442), .I3(rd_addr_r_c[2]), .O(n13769));
    defparam rd_addr_r_1__bdd_4_lut_11735.LUT_INIT = 16'he4aa;
    SB_LUT4 n13067_bdd_4_lut (.I0(n13067), .I1(n11517), .I2(n11516), .I3(rd_addr_r_c[2]), 
            .O(n13070));
    defparam n13067_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i3326_3327 (.Q(\REG.mem_34_8 ), .C(FIFO_CLK_c), .D(n5483));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3323_3324 (.Q(\REG.mem_34_7 ), .C(FIFO_CLK_c), .D(n5482));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3320_3321 (.Q(\REG.mem_34_6 ), .C(FIFO_CLK_c), .D(n5481));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3317_3318 (.Q(\REG.mem_34_5 ), .C(FIFO_CLK_c), .D(n5480));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3314_3315 (.Q(\REG.mem_34_4 ), .C(FIFO_CLK_c), .D(n5479));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3311_3312 (.Q(\REG.mem_34_3 ), .C(FIFO_CLK_c), .D(n5478));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3308_3309 (.Q(\REG.mem_34_2 ), .C(FIFO_CLK_c), .D(n5477));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3305_3306 (.Q(\REG.mem_34_1 ), .C(FIFO_CLK_c), .D(n5476));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3302_3303 (.Q(\REG.mem_34_0 ), .C(FIFO_CLK_c), .D(n5474));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3251_3252 (.Q(\REG.mem_33_15 ), .C(FIFO_CLK_c), .D(n5473));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3248_3249 (.Q(\REG.mem_33_14 ), .C(FIFO_CLK_c), .D(n5472));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3245_3246 (.Q(\REG.mem_33_13 ), .C(FIFO_CLK_c), .D(n5471));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3242_3243 (.Q(\REG.mem_33_12 ), .C(FIFO_CLK_c), .D(n5470));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3239_3240 (.Q(\REG.mem_33_11 ), .C(FIFO_CLK_c), .D(n5469));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3236_3237 (.Q(\REG.mem_33_10 ), .C(FIFO_CLK_c), .D(n5468));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4037_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_30_10 ), .O(n5420));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4037_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13769_bdd_4_lut (.I0(n13769), .I1(n11394), .I2(n11393), .I3(rd_addr_r_c[2]), 
            .O(n12020));
    defparam n13769_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4036_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_30_9 ), .O(n5419));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4036_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11095 (.I0(rd_addr_r_c[1]), .I1(n11429), 
            .I2(n11430), .I3(rd_addr_r_c[2]), .O(n13061));
    defparam rd_addr_r_1__bdd_4_lut_11095.LUT_INIT = 16'he4aa;
    SB_LUT4 i4035_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_30_8 ), .O(n5418));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4035_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11685 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_3 ), 
            .I2(\REG.mem_7_3 ), .I3(rd_addr_r_c[1]), .O(n13763));
    defparam rd_addr_r_0__bdd_4_lut_11685.LUT_INIT = 16'he4aa;
    SB_LUT4 n13763_bdd_4_lut (.I0(n13763), .I1(\REG.mem_5_3 ), .I2(\REG.mem_4_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11041));
    defparam n13763_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i3233_3234 (.Q(\REG.mem_33_9 ), .C(FIFO_CLK_c), .D(n5467));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3230_3231 (.Q(\REG.mem_33_8 ), .C(FIFO_CLK_c), .D(n5466));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3227_3228 (.Q(\REG.mem_33_7 ), .C(FIFO_CLK_c), .D(n5465));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3224_3225 (.Q(\REG.mem_33_6 ), .C(FIFO_CLK_c), .D(n5464));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3221_3222 (.Q(\REG.mem_33_5 ), .C(FIFO_CLK_c), .D(n5463));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3218_3219 (.Q(\REG.mem_33_4 ), .C(FIFO_CLK_c), .D(n5462));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3215_3216 (.Q(\REG.mem_33_3 ), .C(FIFO_CLK_c), .D(n5461));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3212_3213 (.Q(\REG.mem_33_2 ), .C(FIFO_CLK_c), .D(n5460));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3209_3210 (.Q(\REG.mem_33_1 ), .C(FIFO_CLK_c), .D(n5459));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3206_3207 (.Q(\REG.mem_33_0 ), .C(FIFO_CLK_c), .D(n5458));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3155_3156 (.Q(\REG.mem_32_15 ), .C(FIFO_CLK_c), .D(n5457));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3152_3153 (.Q(\REG.mem_32_14 ), .C(FIFO_CLK_c), .D(n5456));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3149_3150 (.Q(\REG.mem_32_13 ), .C(FIFO_CLK_c), .D(n5455));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3146_3147 (.Q(\REG.mem_32_12 ), .C(FIFO_CLK_c), .D(n5454));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3143_3144 (.Q(\REG.mem_32_11 ), .C(FIFO_CLK_c), .D(n5453));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13061_bdd_4_lut (.I0(n13061), .I1(n11412), .I2(n11411), .I3(rd_addr_r_c[2]), 
            .O(n13064));
    defparam n13061_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4034_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_30_7 ), .O(n5417));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4034_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11090 (.I0(rd_addr_r_c[1]), .I1(n11285), 
            .I2(n11286), .I3(rd_addr_r_c[2]), .O(n13055));
    defparam rd_addr_r_1__bdd_4_lut_11090.LUT_INIT = 16'he4aa;
    SB_DFF i3140_3141 (.Q(\REG.mem_32_10 ), .C(FIFO_CLK_c), .D(n5452));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4033_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_30_6 ), .O(n5416));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4033_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3137_3138 (.Q(\REG.mem_32_9 ), .C(FIFO_CLK_c), .D(n5451));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3134_3135 (.Q(\REG.mem_32_8 ), .C(FIFO_CLK_c), .D(n5450));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3131_3132 (.Q(\REG.mem_32_7 ), .C(FIFO_CLK_c), .D(n5449));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3128_3129 (.Q(\REG.mem_32_6 ), .C(FIFO_CLK_c), .D(n5448));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3125_3126 (.Q(\REG.mem_32_5 ), .C(FIFO_CLK_c), .D(n5447));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3122_3123 (.Q(\REG.mem_32_4 ), .C(FIFO_CLK_c), .D(n5446));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3119_3120 (.Q(\REG.mem_32_3 ), .C(FIFO_CLK_c), .D(n5445));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3116_3117 (.Q(\REG.mem_32_2 ), .C(FIFO_CLK_c), .D(n5444));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3113_3114 (.Q(\REG.mem_32_1 ), .C(FIFO_CLK_c), .D(n5443));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3110_3111 (.Q(\REG.mem_32_0 ), .C(FIFO_CLK_c), .D(n5442));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3059_3060 (.Q(\REG.mem_31_15 ), .C(FIFO_CLK_c), .D(n5441));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3056_3057 (.Q(\REG.mem_31_14 ), .C(FIFO_CLK_c), .D(n5440));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3053_3054 (.Q(\REG.mem_31_13 ), .C(FIFO_CLK_c), .D(n5439));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3050_3051 (.Q(\REG.mem_31_12 ), .C(FIFO_CLK_c), .D(n5438));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3047_3048 (.Q(\REG.mem_31_11 ), .C(FIFO_CLK_c), .D(n5437));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11675 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_1 ), 
            .I2(\REG.mem_27_1 ), .I3(rd_addr_r_c[1]), .O(n13757));
    defparam rd_addr_r_0__bdd_4_lut_11675.LUT_INIT = 16'he4aa;
    SB_LUT4 n13757_bdd_4_lut (.I0(n13757), .I1(\REG.mem_25_1 ), .I2(\REG.mem_24_1 ), 
            .I3(rd_addr_r_c[1]), .O(n11455));
    defparam n13757_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13055_bdd_4_lut (.I0(n13055), .I1(n11283), .I2(n11282), .I3(rd_addr_r_c[2]), 
            .O(n13058));
    defparam n13055_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i3044_3045 (.Q(\REG.mem_31_10 ), .C(FIFO_CLK_c), .D(n5436));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4032_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_30_5 ), .O(n5415));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4032_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4031_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_30_4 ), .O(n5414));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4031_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i84_2_lut_3_lut (.I0(n36), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n58));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i84_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11085 (.I0(rd_addr_r_c[1]), .I1(n11489), 
            .I2(n11490), .I3(rd_addr_r_c[2]), .O(n13049));
    defparam rd_addr_r_1__bdd_4_lut_11085.LUT_INIT = 16'he4aa;
    SB_LUT4 i4030_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_30_3 ), .O(n5413));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4030_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3041_3042 (.Q(\REG.mem_31_9 ), .C(FIFO_CLK_c), .D(n5435));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3038_3039 (.Q(\REG.mem_31_8 ), .C(FIFO_CLK_c), .D(n5434));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3035_3036 (.Q(\REG.mem_31_7 ), .C(FIFO_CLK_c), .D(n5433));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3032_3033 (.Q(\REG.mem_31_6 ), .C(FIFO_CLK_c), .D(n5432));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3029_3030 (.Q(\REG.mem_31_5 ), .C(FIFO_CLK_c), .D(n5431));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3026_3027 (.Q(\REG.mem_31_4 ), .C(FIFO_CLK_c), .D(n5430));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3023_3024 (.Q(\REG.mem_31_3 ), .C(FIFO_CLK_c), .D(n5429));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3020_3021 (.Q(\REG.mem_31_2 ), .C(FIFO_CLK_c), .D(n5428));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3017_3018 (.Q(\REG.mem_31_1 ), .C(FIFO_CLK_c), .D(n5427));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3014_3015 (.Q(\REG.mem_31_0 ), .C(FIFO_CLK_c), .D(n5426));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2963_2964 (.Q(\REG.mem_30_15 ), .C(FIFO_CLK_c), .D(n5425));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2960_2961 (.Q(\REG.mem_30_14 ), .C(FIFO_CLK_c), .D(n5424));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2957_2958 (.Q(\REG.mem_30_13 ), .C(FIFO_CLK_c), .D(n5423));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2954_2955 (.Q(\REG.mem_30_12 ), .C(FIFO_CLK_c), .D(n5422));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2951_2952 (.Q(\REG.mem_30_11 ), .C(FIFO_CLK_c), .D(n5421));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2948_2949 (.Q(\REG.mem_30_10 ), .C(FIFO_CLK_c), .D(n5420));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10044_3_lut (.I0(\REG.mem_48_15 ), .I1(\REG.mem_49_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11882));
    defparam i10044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10045_3_lut (.I0(\REG.mem_50_15 ), .I1(\REG.mem_51_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11883));
    defparam i10045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10057_3_lut (.I0(\REG.mem_54_15 ), .I1(\REG.mem_55_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11895));
    defparam i10057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_inv_0_i7_1_lut (.I0(rp_sync2_r[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_45[6]));   // src/fifo_dc_32_lut_gen.v(212[47:78])
    defparam wr_addr_r_6__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4029_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_30_2 ), .O(n5412));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4029_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13049_bdd_4_lut (.I0(n13049), .I1(n11478), .I2(n11477), .I3(rd_addr_r_c[2]), 
            .O(n13052));
    defparam n13049_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10056_3_lut (.I0(\REG.mem_52_15 ), .I1(\REG.mem_53_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11894));
    defparam i10056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4028_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_30_1 ), .O(n5411));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4028_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11670 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_2 ), 
            .I2(\REG.mem_47_2 ), .I3(rd_addr_r_c[1]), .O(n13751));
    defparam rd_addr_r_0__bdd_4_lut_11670.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11080 (.I0(rd_addr_r_c[1]), .I1(n11450), 
            .I2(n11451), .I3(rd_addr_r_c[2]), .O(n13043));
    defparam rd_addr_r_1__bdd_4_lut_11080.LUT_INIT = 16'he4aa;
    SB_DFF i2945_2946 (.Q(\REG.mem_30_9 ), .C(FIFO_CLK_c), .D(n5419));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2942_2943 (.Q(\REG.mem_30_8 ), .C(FIFO_CLK_c), .D(n5418));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2939_2940 (.Q(\REG.mem_30_7 ), .C(FIFO_CLK_c), .D(n5417));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2936_2937 (.Q(\REG.mem_30_6 ), .C(FIFO_CLK_c), .D(n5416));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2933_2934 (.Q(\REG.mem_30_5 ), .C(FIFO_CLK_c), .D(n5415));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2930_2931 (.Q(\REG.mem_30_4 ), .C(FIFO_CLK_c), .D(n5414));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2927_2928 (.Q(\REG.mem_30_3 ), .C(FIFO_CLK_c), .D(n5413));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2924_2925 (.Q(\REG.mem_30_2 ), .C(FIFO_CLK_c), .D(n5412));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2921_2922 (.Q(\REG.mem_30_1 ), .C(FIFO_CLK_c), .D(n5411));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2918_2919 (.Q(\REG.mem_30_0 ), .C(FIFO_CLK_c), .D(n5410));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2867_2868 (.Q(\REG.mem_29_15 ), .C(FIFO_CLK_c), .D(n5409));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2864_2865 (.Q(\REG.mem_29_14 ), .C(FIFO_CLK_c), .D(n5408));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2861_2862 (.Q(\REG.mem_29_13 ), .C(FIFO_CLK_c), .D(n5407));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2858_2859 (.Q(\REG.mem_29_12 ), .C(FIFO_CLK_c), .D(n5406));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2855_2856 (.Q(\REG.mem_29_11 ), .C(FIFO_CLK_c), .D(n5405));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2852_2853 (.Q(\REG.mem_29_10 ), .C(FIFO_CLK_c), .D(n5404));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13043_bdd_4_lut (.I0(n13043), .I1(n11448), .I2(n11447), .I3(rd_addr_r_c[2]), 
            .O(n13046));
    defparam n13043_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4027_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_30_0 ), .O(n5410));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4027_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13751_bdd_4_lut (.I0(n13751), .I1(\REG.mem_45_2 ), .I2(\REG.mem_44_2 ), 
            .I3(rd_addr_r_c[1]), .O(n13754));
    defparam n13751_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4074_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_32_15 ), .O(n5457));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4074_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4073_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_32_14 ), .O(n5456));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4073_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4072_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_32_13 ), .O(n5455));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4072_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11075 (.I0(rd_addr_r_c[1]), .I1(n11243), 
            .I2(n11244), .I3(rd_addr_r_c[2]), .O(n13037));
    defparam rd_addr_r_1__bdd_4_lut_11075.LUT_INIT = 16'he4aa;
    SB_LUT4 i4071_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_32_12 ), .O(n5454));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4071_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4070_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_32_11 ), .O(n5453));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4070_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4069_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_32_10 ), .O(n5452));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4069_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4068_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_32_9 ), .O(n5451));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4068_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11705 (.I0(rd_addr_r_c[3]), .I1(n11921), 
            .I2(n11922), .I3(rd_addr_r_c[4]), .O(n13745));
    defparam rd_addr_r_3__bdd_4_lut_11705.LUT_INIT = 16'he4aa;
    SB_LUT4 n13745_bdd_4_lut (.I0(n13745), .I1(n11901), .I2(n11900), .I3(rd_addr_r_c[4]), 
            .O(n13748));
    defparam n13745_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4067_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_32_8 ), .O(n5450));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4067_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4066_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_32_7 ), .O(n5449));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4066_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4065_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_32_6 ), .O(n5448));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4065_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4064_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_32_5 ), .O(n5447));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4064_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2849_2850 (.Q(\REG.mem_29_9 ), .C(FIFO_CLK_c), .D(n5403));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2846_2847 (.Q(\REG.mem_29_8 ), .C(FIFO_CLK_c), .D(n5402));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2843_2844 (.Q(\REG.mem_29_7 ), .C(FIFO_CLK_c), .D(n5401));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2840_2841 (.Q(\REG.mem_29_6 ), .C(FIFO_CLK_c), .D(n5400));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2837_2838 (.Q(\REG.mem_29_5 ), .C(FIFO_CLK_c), .D(n5399));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2834_2835 (.Q(\REG.mem_29_4 ), .C(FIFO_CLK_c), .D(n5398));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2831_2832 (.Q(\REG.mem_29_3 ), .C(FIFO_CLK_c), .D(n5397));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2828_2829 (.Q(\REG.mem_29_2 ), .C(FIFO_CLK_c), .D(n5396));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2825_2826 (.Q(\REG.mem_29_1 ), .C(FIFO_CLK_c), .D(n5395));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2822_2823 (.Q(\REG.mem_29_0 ), .C(FIFO_CLK_c), .D(n5394));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2771_2772 (.Q(\REG.mem_28_15 ), .C(FIFO_CLK_c), .D(n5393));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2768_2769 (.Q(\REG.mem_28_14 ), .C(FIFO_CLK_c), .D(n5392));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2765_2766 (.Q(\REG.mem_28_13 ), .C(FIFO_CLK_c), .D(n5391));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2762_2763 (.Q(\REG.mem_28_12 ), .C(FIFO_CLK_c), .D(n5390));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2759_2760 (.Q(\REG.mem_28_11 ), .C(FIFO_CLK_c), .D(n5389));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2756_2757 (.Q(\REG.mem_28_10 ), .C(FIFO_CLK_c), .D(n5388));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2753_2754 (.Q(\REG.mem_28_9 ), .C(FIFO_CLK_c), .D(n5387));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13037_bdd_4_lut (.I0(n13037), .I1(n11202), .I2(n11201), .I3(rd_addr_r_c[2]), 
            .O(n13040));
    defparam n13037_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4063_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_32_4 ), .O(n5446));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4063_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4062_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_32_3 ), .O(n5445));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4062_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11665 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_6 ), 
            .I2(\REG.mem_43_6 ), .I3(rd_addr_r_c[1]), .O(n13739));
    defparam rd_addr_r_0__bdd_4_lut_11665.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i83_2_lut_3_lut (.I0(n36), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n26));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i83_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i4061_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_32_2 ), .O(n5444));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4061_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2750_2751 (.Q(\REG.mem_28_8 ), .C(FIFO_CLK_c), .D(n5386));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4060_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_32_1 ), .O(n5443));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4060_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4059_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_32_0 ), .O(n5442));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4059_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13739_bdd_4_lut (.I0(n13739), .I1(\REG.mem_41_6 ), .I2(\REG.mem_40_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11464));
    defparam n13739_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4622_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_62_15 ), .O(n6005));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4622_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11740 (.I0(rd_addr_r_c[2]), .I1(n12938), 
            .I2(n12812), .I3(rd_addr_r_c[3]), .O(n13733));
    defparam rd_addr_r_2__bdd_4_lut_11740.LUT_INIT = 16'he4aa;
    SB_DFF i2747_2748 (.Q(\REG.mem_28_7 ), .C(FIFO_CLK_c), .D(n5385));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2744_2745 (.Q(\REG.mem_28_6 ), .C(FIFO_CLK_c), .D(n5384));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2741_2742 (.Q(\REG.mem_28_5 ), .C(FIFO_CLK_c), .D(n5383));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2738_2739 (.Q(\REG.mem_28_4 ), .C(FIFO_CLK_c), .D(n5382));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2735_2736 (.Q(\REG.mem_28_3 ), .C(FIFO_CLK_c), .D(n5381));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2732_2733 (.Q(\REG.mem_28_2 ), .C(FIFO_CLK_c), .D(n5380));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2729_2730 (.Q(\REG.mem_28_1 ), .C(FIFO_CLK_c), .D(n5379));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2726_2727 (.Q(\REG.mem_28_0 ), .C(FIFO_CLK_c), .D(n5378));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2675_2676 (.Q(\REG.mem_27_15 ), .C(FIFO_CLK_c), .D(n5377));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2672_2673 (.Q(\REG.mem_27_14 ), .C(FIFO_CLK_c), .D(n5376));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2669_2670 (.Q(\REG.mem_27_13 ), .C(FIFO_CLK_c), .D(n5375));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2666_2667 (.Q(\REG.mem_27_12 ), .C(FIFO_CLK_c), .D(n5374));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2663_2664 (.Q(\REG.mem_27_11 ), .C(FIFO_CLK_c), .D(n5373));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2660_2661 (.Q(\REG.mem_27_10 ), .C(FIFO_CLK_c), .D(n5372));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2657_2658 (.Q(\REG.mem_27_9 ), .C(FIFO_CLK_c), .D(n5371));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2654_2655 (.Q(\REG.mem_27_8 ), .C(FIFO_CLK_c), .D(n5370));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i134_135 (.Q(\REG.mem_1_0 ), .C(FIFO_CLK_c), .D(n4884));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11070 (.I0(rd_addr_r_c[1]), .I1(n11423), 
            .I2(n11424), .I3(rd_addr_r_c[2]), .O(n13031));
    defparam rd_addr_r_1__bdd_4_lut_11070.LUT_INIT = 16'he4aa;
    SB_LUT4 i4621_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_62_14 ), .O(n6004));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4621_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13733_bdd_4_lut (.I0(n13733), .I1(n13112), .I2(n13214), .I3(rd_addr_r_c[3]), 
            .O(n11941));
    defparam n13733_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13031_bdd_4_lut (.I0(n13031), .I1(n11415), .I2(n11414), .I3(rd_addr_r_c[2]), 
            .O(n13034));
    defparam n13031_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4620_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_62_13 ), .O(n6003));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4620_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11655 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_0 ), 
            .I2(\REG.mem_47_0 ), .I3(rd_addr_r_c[1]), .O(n13727));
    defparam rd_addr_r_0__bdd_4_lut_11655.LUT_INIT = 16'he4aa;
    SB_DFF i2651_2652 (.Q(\REG.mem_27_7 ), .C(FIFO_CLK_c), .D(n5369));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2648_2649 (.Q(\REG.mem_27_6 ), .C(FIFO_CLK_c), .D(n5368));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2645_2646 (.Q(\REG.mem_27_5 ), .C(FIFO_CLK_c), .D(n5367));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2642_2643 (.Q(\REG.mem_27_4 ), .C(FIFO_CLK_c), .D(n5366));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2639_2640 (.Q(\REG.mem_27_3 ), .C(FIFO_CLK_c), .D(n5365));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2636_2637 (.Q(\REG.mem_27_2 ), .C(FIFO_CLK_c), .D(n5364));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2633_2634 (.Q(\REG.mem_27_1 ), .C(FIFO_CLK_c), .D(n5363));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2630_2631 (.Q(\REG.mem_27_0 ), .C(FIFO_CLK_c), .D(n5362));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2579_2580 (.Q(\REG.mem_26_15 ), .C(FIFO_CLK_c), .D(n5361));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2576_2577 (.Q(\REG.mem_26_14 ), .C(FIFO_CLK_c), .D(n5360));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2573_2574 (.Q(\REG.mem_26_13 ), .C(FIFO_CLK_c), .D(n5359));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2570_2571 (.Q(\REG.mem_26_12 ), .C(FIFO_CLK_c), .D(n5358));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2567_2568 (.Q(\REG.mem_26_11 ), .C(FIFO_CLK_c), .D(n5357));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2564_2565 (.Q(\REG.mem_26_10 ), .C(FIFO_CLK_c), .D(n5356));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2561_2562 (.Q(\REG.mem_26_9 ), .C(FIFO_CLK_c), .D(n5355));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2558_2559 (.Q(\REG.mem_26_8 ), .C(FIFO_CLK_c), .D(n5354));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2555_2556 (.Q(\REG.mem_26_7 ), .C(FIFO_CLK_c), .D(n5353));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4619_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_62_12 ), .O(n6002));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4619_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2552_2553 (.Q(\REG.mem_26_6 ), .C(FIFO_CLK_c), .D(n5352));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4618_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_62_11 ), .O(n6001));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4618_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4617_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_62_10 ), .O(n6000));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4617_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13727_bdd_4_lut (.I0(n13727), .I1(\REG.mem_45_0 ), .I2(\REG.mem_44_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11947));
    defparam n13727_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut (.I0(dc32_fifo_almost_full), .I1(DEBUG_1_c_c), .I2(GND_net), 
            .I3(GND_net), .O(write_to_dc32_fifo_latched_N_425));   // src/fifo_dc_32_lut_gen.v(410[29] 422[32])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11105 (.I0(rd_addr_r_c[3]), .I1(n13010), 
            .I2(n11472), .I3(rd_addr_r_c[4]), .O(n13025));
    defparam rd_addr_r_3__bdd_4_lut_11105.LUT_INIT = 16'he4aa;
    SB_DFF i2549_2550 (.Q(\REG.mem_26_5 ), .C(FIFO_CLK_c), .D(n5351));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4616_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_62_9 ), .O(n5999));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4616_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2546_2547 (.Q(\REG.mem_26_4 ), .C(FIFO_CLK_c), .D(n5350));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2543_2544 (.Q(\REG.mem_26_3 ), .C(FIFO_CLK_c), .D(n5349));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2540_2541 (.Q(\REG.mem_26_2 ), .C(FIFO_CLK_c), .D(n5348));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2537_2538 (.Q(\REG.mem_26_1 ), .C(FIFO_CLK_c), .D(n5347));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2534_2535 (.Q(\REG.mem_26_0 ), .C(FIFO_CLK_c), .D(n5346));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2483_2484 (.Q(\REG.mem_25_15 ), .C(FIFO_CLK_c), .D(n5345));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2480_2481 (.Q(\REG.mem_25_14 ), .C(FIFO_CLK_c), .D(n5344));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2477_2478 (.Q(\REG.mem_25_13 ), .C(FIFO_CLK_c), .D(n5343));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2474_2475 (.Q(\REG.mem_25_12 ), .C(FIFO_CLK_c), .D(n5342));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2471_2472 (.Q(\REG.mem_25_11 ), .C(FIFO_CLK_c), .D(n5341));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2468_2469 (.Q(\REG.mem_25_10 ), .C(FIFO_CLK_c), .D(n5340));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2465_2466 (.Q(\REG.mem_25_9 ), .C(FIFO_CLK_c), .D(n5339));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2462_2463 (.Q(\REG.mem_25_8 ), .C(FIFO_CLK_c), .D(n5338));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2459_2460 (.Q(\REG.mem_25_7 ), .C(FIFO_CLK_c), .D(n5337));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2456_2457 (.Q(\REG.mem_25_6 ), .C(FIFO_CLK_c), .D(n5336));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2453_2454 (.Q(\REG.mem_25_5 ), .C(FIFO_CLK_c), .D(n5335));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12341_bdd_4_lut (.I0(n12341), .I1(\REG.mem_45_5 ), .I2(\REG.mem_44_5 ), 
            .I3(rd_addr_r_c[1]), .O(n12344));
    defparam n12341_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4615_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_62_8 ), .O(n5998));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4615_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4614_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_62_7 ), .O(n5997));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4614_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11645 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_2 ), 
            .I2(\REG.mem_59_2 ), .I3(rd_addr_r_c[1]), .O(n13721));
    defparam rd_addr_r_0__bdd_4_lut_11645.LUT_INIT = 16'he4aa;
    SB_LUT4 n13025_bdd_4_lut (.I0(n13025), .I1(n11460), .I2(n12986), .I3(rd_addr_r_c[4]), 
            .O(n13028));
    defparam n13025_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i1_1_lut (.I0(rd_addr_r[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_DFF i2450_2451 (.Q(\REG.mem_25_4 ), .C(FIFO_CLK_c), .D(n5334));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2447_2448 (.Q(\REG.mem_25_3 ), .C(FIFO_CLK_c), .D(n5333));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i2_1_lut (.I0(rd_addr_r_c[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4613_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_62_6 ), .O(n5996));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4613_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13721_bdd_4_lut (.I0(n13721), .I1(\REG.mem_57_2 ), .I2(\REG.mem_56_2 ), 
            .I3(rd_addr_r_c[1]), .O(n13724));
    defparam n13721_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11065 (.I0(rd_addr_r_c[1]), .I1(n11402), 
            .I2(n11403), .I3(rd_addr_r_c[2]), .O(n13019));
    defparam rd_addr_r_1__bdd_4_lut_11065.LUT_INIT = 16'he4aa;
    SB_LUT4 i4612_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_62_5 ), .O(n5995));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4612_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13019_bdd_4_lut (.I0(n13019), .I1(n11385), .I2(n11384), .I3(rd_addr_r_c[2]), 
            .O(n13022));
    defparam n13019_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i2444_2445 (.Q(\REG.mem_25_2 ), .C(FIFO_CLK_c), .D(n5332));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4611_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_62_4 ), .O(n5994));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4611_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2441_2442 (.Q(\REG.mem_25_1 ), .C(FIFO_CLK_c), .D(n5331));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2438_2439 (.Q(\REG.mem_25_0 ), .C(FIFO_CLK_c), .D(n5330));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10113_3_lut (.I0(n13274), .I1(n13190), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11951));
    defparam i10113_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2387_2388 (.Q(\REG.mem_24_15 ), .C(FIFO_CLK_c), .D(n5329));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2384_2385 (.Q(\REG.mem_24_14 ), .C(FIFO_CLK_c), .D(n5328));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2381_2382 (.Q(\REG.mem_24_13 ), .C(FIFO_CLK_c), .D(n5327));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2378_2379 (.Q(\REG.mem_24_12 ), .C(FIFO_CLK_c), .D(n5326));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2375_2376 (.Q(\REG.mem_24_11 ), .C(FIFO_CLK_c), .D(n5325));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2372_2373 (.Q(\REG.mem_24_10 ), .C(FIFO_CLK_c), .D(n5324));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2369_2370 (.Q(\REG.mem_24_9 ), .C(FIFO_CLK_c), .D(n5323));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2366_2367 (.Q(\REG.mem_24_8 ), .C(FIFO_CLK_c), .D(n5322));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2363_2364 (.Q(\REG.mem_24_7 ), .C(FIFO_CLK_c), .D(n5321));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2360_2361 (.Q(\REG.mem_24_6 ), .C(FIFO_CLK_c), .D(n5320));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2357_2358 (.Q(\REG.mem_24_5 ), .C(FIFO_CLK_c), .D(n5319));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2354_2355 (.Q(\REG.mem_24_4 ), .C(FIFO_CLK_c), .D(n5318));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2351_2352 (.Q(\REG.mem_24_3 ), .C(FIFO_CLK_c), .D(n5317));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2348_2349 (.Q(\REG.mem_24_2 ), .C(FIFO_CLK_c), .D(n5316));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2345_2346 (.Q(\REG.mem_24_1 ), .C(FIFO_CLK_c), .D(n5315));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4610_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_62_3 ), .O(n5993));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4610_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11120 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_15 ), 
            .I2(\REG.mem_15_15 ), .I3(rd_addr_r_c[1]), .O(n13013));
    defparam rd_addr_r_0__bdd_4_lut_11120.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11640 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_13 ), 
            .I2(\REG.mem_7_13 ), .I3(rd_addr_r_c[1]), .O(n13715));
    defparam rd_addr_r_0__bdd_4_lut_11640.LUT_INIT = 16'he4aa;
    SB_LUT4 i4609_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_62_2 ), .O(n5992));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4609_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4608_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_62_1 ), .O(n5991));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4608_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10114_3_lut (.I0(n13136), .I1(n13016), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11952));
    defparam i10114_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2342_2343 (.Q(\REG.mem_24_0 ), .C(FIFO_CLK_c), .D(n5307));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2291_2292 (.Q(\REG.mem_23_15 ), .C(FIFO_CLK_c), .D(n5306));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2288_2289 (.Q(\REG.mem_23_14 ), .C(FIFO_CLK_c), .D(n5305));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2285_2286 (.Q(\REG.mem_23_13 ), .C(FIFO_CLK_c), .D(n5304));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2282_2283 (.Q(\REG.mem_23_12 ), .C(FIFO_CLK_c), .D(n5303));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2279_2280 (.Q(\REG.mem_23_11 ), .C(FIFO_CLK_c), .D(n5302));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2276_2277 (.Q(\REG.mem_23_10 ), .C(FIFO_CLK_c), .D(n5301));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2273_2274 (.Q(\REG.mem_23_9 ), .C(FIFO_CLK_c), .D(n5300));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2270_2271 (.Q(\REG.mem_23_8 ), .C(FIFO_CLK_c), .D(n5299));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2267_2268 (.Q(\REG.mem_23_7 ), .C(FIFO_CLK_c), .D(n5298));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2264_2265 (.Q(\REG.mem_23_6 ), .C(FIFO_CLK_c), .D(n5297));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2261_2262 (.Q(\REG.mem_23_5 ), .C(FIFO_CLK_c), .D(n5296));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2258_2259 (.Q(\REG.mem_23_4 ), .C(FIFO_CLK_c), .D(n5295));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2255_2256 (.Q(\REG.mem_23_3 ), .C(FIFO_CLK_c), .D(n5294));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2252_2253 (.Q(\REG.mem_23_2 ), .C(FIFO_CLK_c), .D(n5293));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2249_2250 (.Q(\REG.mem_23_1 ), .C(FIFO_CLK_c), .D(n5292));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2246_2247 (.Q(\REG.mem_23_0 ), .C(FIFO_CLK_c), .D(n5290));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2195_2196 (.Q(\REG.mem_22_15 ), .C(FIFO_CLK_c), .D(n5289));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2192_2193 (.Q(\REG.mem_22_14 ), .C(FIFO_CLK_c), .D(n5288));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2189_2190 (.Q(\REG.mem_22_13 ), .C(FIFO_CLK_c), .D(n5287));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2186_2187 (.Q(\REG.mem_22_12 ), .C(FIFO_CLK_c), .D(n5286));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2183_2184 (.Q(\REG.mem_22_11 ), .C(FIFO_CLK_c), .D(n5285));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4607_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_62_0 ), .O(n5990));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4607_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFSR rd_grey_sync_r__i5 (.Q(\rd_grey_sync_r[5] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[5]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_LUT4 n13715_bdd_4_lut (.I0(n13715), .I1(\REG.mem_5_13 ), .I2(\REG.mem_4_13 ), 
            .I3(rd_addr_r_c[1]), .O(n11959));
    defparam n13715_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR rd_grey_sync_r__i4 (.Q(\rd_grey_sync_r[4] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[4]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i3 (.Q(\rd_grey_sync_r[3] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[3]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i2 (.Q(\rd_grey_sync_r[2] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[2]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i1 (.Q(\rd_grey_sync_r[1] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[1]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFF i2180_2181 (.Q(\REG.mem_22_10 ), .C(FIFO_CLK_c), .D(n5284));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2177_2178 (.Q(\REG.mem_22_9 ), .C(FIFO_CLK_c), .D(n5283));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2174_2175 (.Q(\REG.mem_22_8 ), .C(FIFO_CLK_c), .D(n5282));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2171_2172 (.Q(\REG.mem_22_7 ), .C(FIFO_CLK_c), .D(n5281));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2168_2169 (.Q(\REG.mem_22_6 ), .C(FIFO_CLK_c), .D(n5280));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2165_2166 (.Q(\REG.mem_22_5 ), .C(FIFO_CLK_c), .D(n5279));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2162_2163 (.Q(\REG.mem_22_4 ), .C(FIFO_CLK_c), .D(n5278));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2159_2160 (.Q(\REG.mem_22_3 ), .C(FIFO_CLK_c), .D(n5277));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2156_2157 (.Q(\REG.mem_22_2 ), .C(FIFO_CLK_c), .D(n5276));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2153_2154 (.Q(\REG.mem_22_1 ), .C(FIFO_CLK_c), .D(n5275));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2150_2151 (.Q(\REG.mem_22_0 ), .C(FIFO_CLK_c), .D(n5274));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2099_2100 (.Q(\REG.mem_21_15 ), .C(FIFO_CLK_c), .D(n5273));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2096_2097 (.Q(\REG.mem_21_14 ), .C(FIFO_CLK_c), .D(n5272));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2093_2094 (.Q(\REG.mem_21_13 ), .C(FIFO_CLK_c), .D(n5271));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2090_2091 (.Q(\REG.mem_21_12 ), .C(FIFO_CLK_c), .D(n5270));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2087_2088 (.Q(\REG.mem_21_11 ), .C(FIFO_CLK_c), .D(n5269));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_4__bdd_4_lut_11725 (.I0(rd_addr_r_c[4]), .I1(n11905), 
            .I2(n11941), .I3(rd_addr_r_c[5]), .O(n13709));
    defparam rd_addr_r_4__bdd_4_lut_11725.LUT_INIT = 16'he4aa;
    SB_LUT4 n13013_bdd_4_lut (.I0(n13013), .I1(\REG.mem_13_15 ), .I2(\REG.mem_12_15 ), 
            .I3(rd_addr_r_c[1]), .O(n13016));
    defparam n13013_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13709_bdd_4_lut (.I0(n13709), .I1(n12290), .I2(n12458), .I3(rd_addr_r_c[5]), 
            .O(\REG.out_raw_31__N_559 [1]));
    defparam n13709_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i98_2_lut_3_lut_4_lut (.I0(n17_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n51));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i98_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_DFF i2084_2085 (.Q(\REG.mem_21_10 ), .C(FIFO_CLK_c), .D(n5268));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2081_2082 (.Q(\REG.mem_21_9 ), .C(FIFO_CLK_c), .D(n5267));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2078_2079 (.Q(\REG.mem_21_8 ), .C(FIFO_CLK_c), .D(n5266));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2075_2076 (.Q(\REG.mem_21_7 ), .C(FIFO_CLK_c), .D(n5265));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2072_2073 (.Q(\REG.mem_21_6 ), .C(FIFO_CLK_c), .D(n5264));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2069_2070 (.Q(\REG.mem_21_5 ), .C(FIFO_CLK_c), .D(n5263));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2066_2067 (.Q(\REG.mem_21_4 ), .C(FIFO_CLK_c), .D(n5262));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2063_2064 (.Q(\REG.mem_21_3 ), .C(FIFO_CLK_c), .D(n5261));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2060_2061 (.Q(\REG.mem_21_2 ), .C(FIFO_CLK_c), .D(n5260));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2057_2058 (.Q(\REG.mem_21_1 ), .C(FIFO_CLK_c), .D(n5259));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2054_2055 (.Q(\REG.mem_21_0 ), .C(FIFO_CLK_c), .D(n5257));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2003_2004 (.Q(\REG.mem_20_15 ), .C(FIFO_CLK_c), .D(n5256));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2000_2001 (.Q(\REG.mem_20_14 ), .C(FIFO_CLK_c), .D(n5255));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1997_1998 (.Q(\REG.mem_20_13 ), .C(FIFO_CLK_c), .D(n5254));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1994_1995 (.Q(\REG.mem_20_12 ), .C(FIFO_CLK_c), .D(n5253));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i97_2_lut_3_lut_4_lut (.I0(n17_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n19));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i97_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i4603_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_61_15 ), .O(n5986));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4603_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4602_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_61_14 ), .O(n5985));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4602_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1991_1992 (.Q(\REG.mem_20_11 ), .C(FIFO_CLK_c), .D(n5252));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11055 (.I0(rd_addr_r_c[1]), .I1(n11204), 
            .I2(n11205), .I3(rd_addr_r_c[2]), .O(n13007));
    defparam rd_addr_r_1__bdd_4_lut_11055.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11635 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_13 ), 
            .I2(\REG.mem_47_13 ), .I3(rd_addr_r_c[1]), .O(n13703));
    defparam rd_addr_r_0__bdd_4_lut_11635.LUT_INIT = 16'he4aa;
    SB_LUT4 n13703_bdd_4_lut (.I0(n13703), .I1(\REG.mem_45_13 ), .I2(\REG.mem_44_13 ), 
            .I3(rd_addr_r_c[1]), .O(n11482));
    defparam n13703_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13007_bdd_4_lut (.I0(n13007), .I1(n11163), .I2(n11162), .I3(rd_addr_r_c[2]), 
            .O(n13010));
    defparam n13007_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11625 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_2 ), 
            .I2(\REG.mem_63_2 ), .I3(rd_addr_r_c[1]), .O(n13697));
    defparam rd_addr_r_0__bdd_4_lut_11625.LUT_INIT = 16'he4aa;
    SB_LUT4 i4601_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_61_13 ), .O(n5984));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4601_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4600_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_61_12 ), .O(n5983));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4600_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13697_bdd_4_lut (.I0(n13697), .I1(\REG.mem_61_2 ), .I2(\REG.mem_60_2 ), 
            .I3(rd_addr_r_c[1]), .O(n13700));
    defparam n13697_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4599_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_61_11 ), .O(n5982));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4599_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4598_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_61_10 ), .O(n5981));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4598_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4597_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_61_9 ), .O(n5980));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4597_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4596_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_61_8 ), .O(n5979));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4596_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1988_1989 (.Q(\REG.mem_20_10 ), .C(FIFO_CLK_c), .D(n5251));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11620 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_6 ), 
            .I2(\REG.mem_47_6 ), .I3(rd_addr_r_c[1]), .O(n13691));
    defparam rd_addr_r_0__bdd_4_lut_11620.LUT_INIT = 16'he4aa;
    SB_DFF i1985_1986 (.Q(\REG.mem_20_9 ), .C(FIFO_CLK_c), .D(n5250));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1982_1983 (.Q(\REG.mem_20_8 ), .C(FIFO_CLK_c), .D(n5249));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1979_1980 (.Q(\REG.mem_20_7 ), .C(FIFO_CLK_c), .D(n5248));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1976_1977 (.Q(\REG.mem_20_6 ), .C(FIFO_CLK_c), .D(n5247));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1973_1974 (.Q(\REG.mem_20_5 ), .C(FIFO_CLK_c), .D(n5246));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1970_1971 (.Q(\REG.mem_20_4 ), .C(FIFO_CLK_c), .D(n5245));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1967_1968 (.Q(\REG.mem_20_3 ), .C(FIFO_CLK_c), .D(n5244));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1964_1965 (.Q(\REG.mem_20_2 ), .C(FIFO_CLK_c), .D(n5243));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1961_1962 (.Q(\REG.mem_20_1 ), .C(FIFO_CLK_c), .D(n5242));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1958_1959 (.Q(\REG.mem_20_0 ), .C(FIFO_CLK_c), .D(n5241));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1907_1908 (.Q(\REG.mem_19_15 ), .C(FIFO_CLK_c), .D(n5240));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1904_1905 (.Q(\REG.mem_19_14 ), .C(FIFO_CLK_c), .D(n5239));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1901_1902 (.Q(\REG.mem_19_13 ), .C(FIFO_CLK_c), .D(n5238));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1898_1899 (.Q(\REG.mem_19_12 ), .C(FIFO_CLK_c), .D(n5237));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4595_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_61_7 ), .O(n5978));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4595_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4594_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_61_6 ), .O(n5977));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4594_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_r_6__I_0_135_i2_3_lut (.I0(wr_addr_r[1]), .I1(wr_addr_p1_w[1]), 
            .I2(wr_sig_mv_w), .I3(GND_net), .O(\wr_addr_nxt_c[1] ));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_6__I_0_135_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11050 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_12 ), 
            .I2(\REG.mem_35_12 ), .I3(rd_addr_r_c[1]), .O(n13001));
    defparam rd_addr_r_0__bdd_4_lut_11050.LUT_INIT = 16'he4aa;
    SB_LUT4 i4593_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_61_5 ), .O(n5976));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4593_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4592_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_61_4 ), .O(n5975));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4592_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13691_bdd_4_lut (.I0(n13691), .I1(\REG.mem_45_6 ), .I2(\REG.mem_44_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11485));
    defparam n13691_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13001_bdd_4_lut (.I0(n13001), .I1(\REG.mem_33_12 ), .I2(\REG.mem_32_12 ), 
            .I3(rd_addr_r_c[1]), .O(n13004));
    defparam n13001_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4591_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_61_3 ), .O(n5974));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4591_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4590_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_61_2 ), .O(n5973));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4590_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4090_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_33_15 ), .O(n5473));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4090_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11040 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_0 ), 
            .I2(\REG.mem_11_0 ), .I3(rd_addr_r_c[1]), .O(n12995));
    defparam rd_addr_r_0__bdd_4_lut_11040.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11615 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_3 ), 
            .I2(\REG.mem_11_3 ), .I3(rd_addr_r_c[1]), .O(n13685));
    defparam rd_addr_r_0__bdd_4_lut_11615.LUT_INIT = 16'he4aa;
    SB_DFF i1895_1896 (.Q(\REG.mem_19_11 ), .C(FIFO_CLK_c), .D(n5236));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4589_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_61_1 ), .O(n5972));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4589_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4588_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_61_0 ), .O(n5971));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4588_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1892_1893 (.Q(\REG.mem_19_10 ), .C(FIFO_CLK_c), .D(n5235));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1889_1890 (.Q(\REG.mem_19_9 ), .C(FIFO_CLK_c), .D(n5234));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1886_1887 (.Q(\REG.mem_19_8 ), .C(FIFO_CLK_c), .D(n5233));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1883_1884 (.Q(\REG.mem_19_7 ), .C(FIFO_CLK_c), .D(n5232));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1880_1881 (.Q(\REG.mem_19_6 ), .C(FIFO_CLK_c), .D(n5231));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1877_1878 (.Q(\REG.mem_19_5 ), .C(FIFO_CLK_c), .D(n5230));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1874_1875 (.Q(\REG.mem_19_4 ), .C(FIFO_CLK_c), .D(n5229));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1871_1872 (.Q(\REG.mem_19_3 ), .C(FIFO_CLK_c), .D(n5228));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1868_1869 (.Q(\REG.mem_19_2 ), .C(FIFO_CLK_c), .D(n5227));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1865_1866 (.Q(\REG.mem_19_1 ), .C(FIFO_CLK_c), .D(n5226));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1862_1863 (.Q(\REG.mem_19_0 ), .C(FIFO_CLK_c), .D(n5225));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1811_1812 (.Q(\REG.mem_18_15 ), .C(FIFO_CLK_c), .D(n5224));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1808_1809 (.Q(\REG.mem_18_14 ), .C(FIFO_CLK_c), .D(n5223));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1805_1806 (.Q(\REG.mem_18_13 ), .C(FIFO_CLK_c), .D(n5222));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1802_1803 (.Q(\REG.mem_18_12 ), .C(FIFO_CLK_c), .D(n5221));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1799_1800 (.Q(\REG.mem_18_11 ), .C(FIFO_CLK_c), .D(n5220));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i1_2_lut_adj_28 (.I0(wp_sync2_r[1]), .I1(wp_sync_w[2]), .I2(GND_net), 
            .I3(GND_net), .O(wp_sync_w[1]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_28.LUT_INIT = 16'h6666;
    SB_LUT4 n13685_bdd_4_lut (.I0(n13685), .I1(\REG.mem_9_3 ), .I2(\REG.mem_8_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11044));
    defparam n13685_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12995_bdd_4_lut (.I0(n12995), .I1(\REG.mem_9_0 ), .I2(\REG.mem_8_0 ), 
            .I3(rd_addr_r_c[1]), .O(n12998));
    defparam n12995_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11610 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_13 ), 
            .I2(\REG.mem_11_13 ), .I3(rd_addr_r_c[1]), .O(n13679));
    defparam rd_addr_r_0__bdd_4_lut_11610.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i96_2_lut_3_lut_4_lut (.I0(n15_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n52));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i96_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 n13679_bdd_4_lut (.I0(n13679), .I1(\REG.mem_9_13 ), .I2(\REG.mem_8_13 ), 
            .I3(rd_addr_r_c[1]), .O(n11965));
    defparam n13679_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i95_2_lut_3_lut_4_lut (.I0(n15_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n20));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i95_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_adj_29 (.I0(wp_sync2_r[3]), .I1(wp_sync_w[4]), .I2(GND_net), 
            .I3(GND_net), .O(wp_sync_w[3]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_29.LUT_INIT = 16'h6666;
    SB_DFF i1796_1797 (.Q(\REG.mem_18_10 ), .C(FIFO_CLK_c), .D(n5219));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i1_2_lut_adj_30 (.I0(wp_sync2_r[6]), .I1(wp_sync2_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n4274));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_30.LUT_INIT = 16'h6666;
    SB_DFF i1793_1794 (.Q(\REG.mem_18_9 ), .C(FIFO_CLK_c), .D(n5218));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1790_1791 (.Q(\REG.mem_18_8 ), .C(FIFO_CLK_c), .D(n5217));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1787_1788 (.Q(\REG.mem_18_7 ), .C(FIFO_CLK_c), .D(n5216));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1784_1785 (.Q(\REG.mem_18_6 ), .C(FIFO_CLK_c), .D(n5215));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1781_1782 (.Q(\REG.mem_18_5 ), .C(FIFO_CLK_c), .D(n5214));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1778_1779 (.Q(\REG.mem_18_4 ), .C(FIFO_CLK_c), .D(n5213));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1775_1776 (.Q(\REG.mem_18_3 ), .C(FIFO_CLK_c), .D(n5212));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1772_1773 (.Q(\REG.mem_18_2 ), .C(FIFO_CLK_c), .D(n5211));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1769_1770 (.Q(\REG.mem_18_1 ), .C(FIFO_CLK_c), .D(n5210));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1766_1767 (.Q(\REG.mem_18_0 ), .C(FIFO_CLK_c), .D(n5209));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1715_1716 (.Q(\REG.mem_17_15 ), .C(FIFO_CLK_c), .D(n5208));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1712_1713 (.Q(\REG.mem_17_14 ), .C(FIFO_CLK_c), .D(n5207));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1709_1710 (.Q(\REG.mem_17_13 ), .C(FIFO_CLK_c), .D(n5206));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1706_1707 (.Q(\REG.mem_17_12 ), .C(FIFO_CLK_c), .D(n5205));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1703_1704 (.Q(\REG.mem_17_11 ), .C(FIFO_CLK_c), .D(n5204));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9053_4_lut (.I0(rd_addr_r[0]), .I1(rd_addr_r_c[4]), .I2(wp_sync_w[0]), 
            .I3(wp_sync_w[4]), .O(n10889));
    defparam i9053_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i9062_4_lut (.I0(rd_addr_r_c[5]), .I1(rd_addr_r_c[3]), .I2(n4274), 
            .I3(wp_sync_w[3]), .O(n10899));
    defparam i9062_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11605 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_0 ), 
            .I2(\REG.mem_51_0 ), .I3(rd_addr_r_c[1]), .O(n13673));
    defparam rd_addr_r_0__bdd_4_lut_11605.LUT_INIT = 16'he4aa;
    SB_LUT4 i3567_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_2_5 ), .O(n4950));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3567_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3566_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_2_4 ), .O(n4949));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3566_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3532_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_1_11 ), .O(n4915));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3532_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1700_1701 (.Q(\REG.mem_17_10 ), .C(FIFO_CLK_c), .D(n5203));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13673_bdd_4_lut (.I0(n13673), .I1(\REG.mem_49_0 ), .I2(\REG.mem_48_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11968));
    defparam n13673_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_31 (.I0(rd_addr_p1_w[4]), .I1(wp_sync_w[4]), .I2(GND_net), 
            .I3(GND_net), .O(n4298));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_31.LUT_INIT = 16'h6666;
    SB_LUT4 i3565_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_2_3 ), .O(n4948));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3565_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3564_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_2_2 ), .O(n4947));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3564_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut (.I0(rd_addr_p1_w[5]), .I1(rd_addr_p1_w[3]), .I2(n4274), 
            .I3(wp_sync_w[3]), .O(n10_c));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i3_4_lut.LUT_INIT = 16'h7bde;
    SB_DFF i1697_1698 (.Q(\REG.mem_17_9 ), .C(FIFO_CLK_c), .D(n5202));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3563_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_2_1 ), .O(n4946));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3563_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11600 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_13 ), 
            .I2(\REG.mem_15_13 ), .I3(rd_addr_r_c[1]), .O(n13667));
    defparam rd_addr_r_0__bdd_4_lut_11600.LUT_INIT = 16'he4aa;
    SB_LUT4 i3562_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_2_0 ), .O(n4945));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3562_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_32 (.I0(wp_sync2_r[6]), .I1(rd_addr_p1_w[1]), .I2(rd_addr_p1_w[6]), 
            .I3(wp_sync_w[1]), .O(n8_adj_25));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i1_4_lut_adj_32.LUT_INIT = 16'h7bde;
    SB_LUT4 i5_4_lut (.I0(\rd_addr_p1_w[0] ), .I1(n10_c), .I2(n4298), 
            .I3(wp_sync_w[0]), .O(n12));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i5_4_lut.LUT_INIT = 16'hfdfe;
    SB_DFF i1694_1695 (.Q(\REG.mem_17_8 ), .C(FIFO_CLK_c), .D(n5201));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9147_3_lut (.I0(n10887), .I1(n10899), .I2(n10889), .I3(GND_net), 
            .O(n10985));
    defparam i9147_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3577_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_2_15 ), .O(n4960));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3577_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13667_bdd_4_lut (.I0(n13667), .I1(\REG.mem_13_13 ), .I2(\REG.mem_12_13 ), 
            .I3(rd_addr_r_c[1]), .O(n11971));
    defparam n13667_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11035 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_9 ), 
            .I2(\REG.mem_43_9 ), .I3(rd_addr_r_c[1]), .O(n12989));
    defparam rd_addr_r_0__bdd_4_lut_11035.LUT_INIT = 16'he4aa;
    SB_LUT4 n12989_bdd_4_lut (.I0(n12989), .I1(\REG.mem_41_9 ), .I2(\REG.mem_40_9 ), 
            .I3(rd_addr_r_c[1]), .O(n12992));
    defparam n12989_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11595 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_4 ), 
            .I2(\REG.mem_7_4 ), .I3(rd_addr_r_c[1]), .O(n13661));
    defparam rd_addr_r_0__bdd_4_lut_11595.LUT_INIT = 16'he4aa;
    SB_LUT4 n13661_bdd_4_lut (.I0(n13661), .I1(\REG.mem_5_4 ), .I2(\REG.mem_4_4 ), 
            .I3(rd_addr_r_c[1]), .O(n13664));
    defparam n13661_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11045 (.I0(rd_addr_r_c[1]), .I1(n11072), 
            .I2(n11073), .I3(rd_addr_r_c[2]), .O(n12983));
    defparam rd_addr_r_1__bdd_4_lut_11045.LUT_INIT = 16'he4aa;
    SB_LUT4 i6_4_lut (.I0(rd_addr_p1_w[2]), .I1(n12), .I2(n8_adj_25), 
            .I3(wp_sync_w[2]), .O(n10258));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i6_4_lut.LUT_INIT = 16'hfdfe;
    SB_LUT4 i3576_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_2_14 ), .O(n4959));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3576_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1691_1692 (.Q(\REG.mem_17_7 ), .C(FIFO_CLK_c), .D(n5200));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1688_1689 (.Q(\REG.mem_17_6 ), .C(FIFO_CLK_c), .D(n5199));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1685_1686 (.Q(\REG.mem_17_5 ), .C(FIFO_CLK_c), .D(n5198));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1682_1683 (.Q(\REG.mem_17_4 ), .C(FIFO_CLK_c), .D(n5197));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1679_1680 (.Q(\REG.mem_17_3 ), .C(FIFO_CLK_c), .D(n5196));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1676_1677 (.Q(\REG.mem_17_2 ), .C(FIFO_CLK_c), .D(n5195));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1673_1674 (.Q(\REG.mem_17_1 ), .C(FIFO_CLK_c), .D(n5194));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 empty_nxt_c_I_7_4_lut (.I0(n10258), .I1(n10985), .I2(DEBUG_3_c), 
            .I3(get_next_word), .O(empty_nxt_c_N_629));   // src/fifo_dc_32_lut_gen.v(555[46:103])
    defparam empty_nxt_c_I_7_4_lut.LUT_INIT = 16'h3530;
    SB_DFF i1670_1671 (.Q(\REG.mem_17_0 ), .C(FIFO_CLK_c), .D(n5193));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1619_1620 (.Q(\REG.mem_16_15 ), .C(FIFO_CLK_c), .D(n5188));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1616_1617 (.Q(\REG.mem_16_14 ), .C(FIFO_CLK_c), .D(n5186));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3575_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_2_13 ), .O(n4958));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3575_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9178_3_lut (.I0(n12740), .I1(n12668), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11016));
    defparam i9178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10173_3_lut (.I0(\REG.mem_0_6 ), .I1(\REG.mem_1_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12011));
    defparam i10173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3574_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_2_12 ), .O(n4957));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3574_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1613_1614 (.Q(\REG.mem_16_13 ), .C(FIFO_CLK_c), .D(n5185));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11590 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_8 ), 
            .I2(\REG.mem_7_8 ), .I3(rd_addr_r_c[1]), .O(n13655));
    defparam rd_addr_r_0__bdd_4_lut_11590.LUT_INIT = 16'he4aa;
    SB_LUT4 i10174_3_lut (.I0(\REG.mem_2_6 ), .I1(\REG.mem_3_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12012));
    defparam i10174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4089_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_33_14 ), .O(n5472));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4089_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1610_1611 (.Q(\REG.mem_16_12 ), .C(FIFO_CLK_c), .D(n5184));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3573_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_2_11 ), .O(n4956));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3573_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13655_bdd_4_lut (.I0(n13655), .I1(\REG.mem_5_8 ), .I2(\REG.mem_4_8 ), 
            .I3(rd_addr_r_c[1]), .O(n13658));
    defparam n13655_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3572_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_2_10 ), .O(n4955));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3572_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10534 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_2 ), 
            .I2(\REG.mem_7_2 ), .I3(rd_addr_r_c[1]), .O(n12383));
    defparam rd_addr_r_0__bdd_4_lut_10534.LUT_INIT = 16'he4aa;
    SB_LUT4 i3571_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_2_9 ), .O(n4954));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3571_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12383_bdd_4_lut (.I0(n12383), .I1(\REG.mem_5_2 ), .I2(\REG.mem_4_2 ), 
            .I3(rd_addr_r_c[1]), .O(n12386));
    defparam n12383_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11680 (.I0(rd_addr_r_c[1]), .I1(n11936), 
            .I2(n11937), .I3(rd_addr_r_c[2]), .O(n13649));
    defparam rd_addr_r_1__bdd_4_lut_11680.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10529 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_9 ), 
            .I2(\REG.mem_63_9 ), .I3(rd_addr_r_c[1]), .O(n12377));
    defparam rd_addr_r_0__bdd_4_lut_10529.LUT_INIT = 16'he4aa;
    SB_LUT4 n12377_bdd_4_lut (.I0(n12377), .I1(\REG.mem_61_9 ), .I2(\REG.mem_60_9 ), 
            .I3(rd_addr_r_c[1]), .O(n12380));
    defparam n12377_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3570_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_2_8 ), .O(n4953));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3570_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3569_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_2_7 ), .O(n4952));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3569_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12983_bdd_4_lut (.I0(n12983), .I1(n11037), .I2(n11036), .I3(rd_addr_r_c[2]), 
            .O(n12986));
    defparam n12983_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13649_bdd_4_lut (.I0(n13649), .I1(n11874), .I2(n11873), .I3(rd_addr_r_c[2]), 
            .O(n11049));
    defparam n13649_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3519_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_1_13 ), .O(n4902));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3519_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3568_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_2_6 ), .O(n4951));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3568_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_6__I_0_i1_3_lut (.I0(rd_addr_r[0]), .I1(\rd_addr_p1_w[0] ), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(rd_addr_nxt_c_6__N_498[0]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_6__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1607_1608 (.Q(\REG.mem_16_11 ), .C(FIFO_CLK_c), .D(n5183));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1604_1605 (.Q(\REG.mem_16_10 ), .C(FIFO_CLK_c), .D(n5182));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1601_1602 (.Q(\REG.mem_16_9 ), .C(FIFO_CLK_c), .D(n5181));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1598_1599 (.Q(\REG.mem_16_8 ), .C(FIFO_CLK_c), .D(n5180));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1595_1596 (.Q(\REG.mem_16_7 ), .C(FIFO_CLK_c), .D(n5179));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1592_1593 (.Q(\REG.mem_16_6 ), .C(FIFO_CLK_c), .D(n5178));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1589_1590 (.Q(\REG.mem_16_5 ), .C(FIFO_CLK_c), .D(n5177));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11585 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_1 ), 
            .I2(\REG.mem_31_1 ), .I3(rd_addr_r_c[1]), .O(n13643));
    defparam rd_addr_r_0__bdd_4_lut_11585.LUT_INIT = 16'he4aa;
    SB_LUT4 n13643_bdd_4_lut (.I0(n13643), .I1(\REG.mem_29_1 ), .I2(\REG.mem_28_1 ), 
            .I3(rd_addr_r_c[1]), .O(n11488));
    defparam n13643_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1586_1587 (.Q(\REG.mem_16_4 ), .C(FIFO_CLK_c), .D(n5176));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i137_138 (.Q(\REG.mem_1_1 ), .C(FIFO_CLK_c), .D(n4879));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4088_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_33_13 ), .O(n5471));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4088_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3529_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_1_12 ), .O(n4912));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3529_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11575 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_13 ), 
            .I2(\REG.mem_51_13 ), .I3(rd_addr_r_c[1]), .O(n13637));
    defparam rd_addr_r_0__bdd_4_lut_11575.LUT_INIT = 16'he4aa;
    SB_LUT4 i10029_3_lut (.I0(\REG.mem_16_14 ), .I1(\REG.mem_17_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11867));
    defparam i10029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10030_3_lut (.I0(\REG.mem_18_14 ), .I1(\REG.mem_19_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11868));
    defparam i10030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9702_3_lut (.I0(\REG.mem_0_12 ), .I1(\REG.mem_1_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11540));
    defparam i9702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13637_bdd_4_lut (.I0(n13637), .I1(\REG.mem_49_13 ), .I2(\REG.mem_48_13 ), 
            .I3(rd_addr_r_c[1]), .O(n11500));
    defparam n13637_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9703_3_lut (.I0(\REG.mem_2_12 ), .I1(\REG.mem_3_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11541));
    defparam i9703_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1583_1584 (.Q(\REG.mem_16_3 ), .C(FIFO_CLK_c), .D(n5175));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1580_1581 (.Q(\REG.mem_16_2 ), .C(FIFO_CLK_c), .D(n5174));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1577_1578 (.Q(\REG.mem_16_1 ), .C(FIFO_CLK_c), .D(n5173));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1574_1575 (.Q(\REG.mem_16_0 ), .C(FIFO_CLK_c), .D(n5172));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1523_1524 (.Q(\REG.mem_15_15 ), .C(FIFO_CLK_c), .D(n5169));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1520_1521 (.Q(\REG.mem_15_14 ), .C(FIFO_CLK_c), .D(n5168));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1517_1518 (.Q(\REG.mem_15_13 ), .C(FIFO_CLK_c), .D(n5167));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i106_2_lut_3_lut_4_lut (.I0(n18_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n47));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i106_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11030 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_11 ), 
            .I2(\REG.mem_43_11 ), .I3(rd_addr_r_c[1]), .O(n12977));
    defparam rd_addr_r_0__bdd_4_lut_11030.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11580 (.I0(rd_addr_r_c[1]), .I1(n11927), 
            .I2(n11928), .I3(rd_addr_r_c[2]), .O(n13631));
    defparam rd_addr_r_1__bdd_4_lut_11580.LUT_INIT = 16'he4aa;
    SB_DFF i1514_1515 (.Q(\REG.mem_15_12 ), .C(FIFO_CLK_c), .D(n5166));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i105_2_lut_3_lut_4_lut (.I0(n18_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n15));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i105_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_DFF i1511_1512 (.Q(\REG.mem_15_11 ), .C(FIFO_CLK_c), .D(n5165));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1508_1509 (.Q(\REG.mem_15_10 ), .C(FIFO_CLK_c), .D(n5164));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1505_1506 (.Q(\REG.mem_15_9 ), .C(FIFO_CLK_c), .D(n5163));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1502_1503 (.Q(\REG.mem_15_8 ), .C(FIFO_CLK_c), .D(n5162));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13631_bdd_4_lut (.I0(n13631), .I1(n11919), .I2(n11918), .I3(rd_addr_r_c[2]), 
            .O(n11052));
    defparam n13631_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1499_1500 (.Q(\REG.mem_15_7 ), .C(FIFO_CLK_c), .D(n5161));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3448_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_1_10 ), .O(n4831));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3448_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12977_bdd_4_lut (.I0(n12977), .I1(\REG.mem_41_11 ), .I2(\REG.mem_40_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11692));
    defparam n12977_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1496_1497 (.Q(\REG.mem_15_6 ), .C(FIFO_CLK_c), .D(n5160));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1493_1494 (.Q(\REG.mem_15_5 ), .C(FIFO_CLK_c), .D(n5159));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1490_1491 (.Q(\REG.mem_15_4 ), .C(FIFO_CLK_c), .D(n5158));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1487_1488 (.Q(\REG.mem_15_3 ), .C(FIFO_CLK_c), .D(n5157));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1484_1485 (.Q(\REG.mem_15_2 ), .C(FIFO_CLK_c), .D(n5156));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1481_1482 (.Q(\REG.mem_15_1 ), .C(FIFO_CLK_c), .D(n5155));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11020 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_12 ), 
            .I2(\REG.mem_39_12 ), .I3(rd_addr_r_c[1]), .O(n12971));
    defparam rd_addr_r_0__bdd_4_lut_11020.LUT_INIT = 16'he4aa;
    SB_DFF i1478_1479 (.Q(\REG.mem_15_0 ), .C(FIFO_CLK_c), .D(n5154));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1427_1428 (.Q(\REG.mem_14_15 ), .C(FIFO_CLK_c), .D(n5153));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1424_1425 (.Q(\REG.mem_14_14 ), .C(FIFO_CLK_c), .D(n5152));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4586_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_60_15 ), .O(n5969));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4586_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4585_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_60_14 ), .O(n5968));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4585_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10186_3_lut (.I0(\REG.mem_6_6 ), .I1(\REG.mem_7_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12024));
    defparam i10186_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1421_1422 (.Q(\REG.mem_14_13 ), .C(FIFO_CLK_c), .D(n5151));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1418_1419 (.Q(\REG.mem_14_12 ), .C(FIFO_CLK_c), .D(n5150));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1415_1416 (.Q(\REG.mem_14_11 ), .C(FIFO_CLK_c), .D(n5149));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1412_1413 (.Q(\REG.mem_14_10 ), .C(FIFO_CLK_c), .D(n5148));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1409_1410 (.Q(\REG.mem_14_9 ), .C(FIFO_CLK_c), .D(n5147));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1406_1407 (.Q(\REG.mem_14_8 ), .C(FIFO_CLK_c), .D(n5146));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1403_1404 (.Q(\REG.mem_14_7 ), .C(FIFO_CLK_c), .D(n5145));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1400_1401 (.Q(\REG.mem_14_6 ), .C(FIFO_CLK_c), .D(n5144));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10185_3_lut (.I0(\REG.mem_4_6 ), .I1(\REG.mem_5_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12023));
    defparam i10185_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1397_1398 (.Q(\REG.mem_14_5 ), .C(FIFO_CLK_c), .D(n5143));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4584_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_60_13 ), .O(n5967));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4584_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1394_1395 (.Q(\REG.mem_14_4 ), .C(FIFO_CLK_c), .D(n5142));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11570 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_9 ), 
            .I2(\REG.mem_15_9 ), .I3(rd_addr_r_c[1]), .O(n13625));
    defparam rd_addr_r_0__bdd_4_lut_11570.LUT_INIT = 16'he4aa;
    SB_DFF i1391_1392 (.Q(\REG.mem_14_3 ), .C(FIFO_CLK_c), .D(n5141));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12971_bdd_4_lut (.I0(n12971), .I1(\REG.mem_37_12 ), .I2(\REG.mem_36_12 ), 
            .I3(rd_addr_r_c[1]), .O(n12974));
    defparam n12971_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1388_1389 (.Q(\REG.mem_14_2 ), .C(FIFO_CLK_c), .D(n5140));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1385_1386 (.Q(\REG.mem_14_1 ), .C(FIFO_CLK_c), .D(n5139));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1382_1383 (.Q(\REG.mem_14_0 ), .C(FIFO_CLK_c), .D(n5138));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1331_1332 (.Q(\REG.mem_13_15 ), .C(FIFO_CLK_c), .D(n5137));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1328_1329 (.Q(\REG.mem_13_14 ), .C(FIFO_CLK_c), .D(n5136));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1325_1326 (.Q(\REG.mem_13_13 ), .C(FIFO_CLK_c), .D(n5135));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1322_1323 (.Q(\REG.mem_13_12 ), .C(FIFO_CLK_c), .D(n5134));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1319_1320 (.Q(\REG.mem_13_11 ), .C(FIFO_CLK_c), .D(n5133));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1316_1317 (.Q(\REG.mem_13_10 ), .C(FIFO_CLK_c), .D(n5132));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13625_bdd_4_lut (.I0(n13625), .I1(\REG.mem_13_9 ), .I2(\REG.mem_12_9 ), 
            .I3(rd_addr_r_c[1]), .O(n11176));
    defparam n13625_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1313_1314 (.Q(\REG.mem_13_9 ), .C(FIFO_CLK_c), .D(n5131));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11560 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_8 ), 
            .I2(\REG.mem_27_8 ), .I3(rd_addr_r_c[1]), .O(n13619));
    defparam rd_addr_r_0__bdd_4_lut_11560.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11015 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_11 ), 
            .I2(\REG.mem_47_11 ), .I3(rd_addr_r_c[1]), .O(n12965));
    defparam rd_addr_r_0__bdd_4_lut_11015.LUT_INIT = 16'he4aa;
    SB_LUT4 n12965_bdd_4_lut (.I0(n12965), .I1(\REG.mem_45_11 ), .I2(\REG.mem_44_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11701));
    defparam n12965_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11025 (.I0(rd_addr_r_c[1]), .I1(n11279), 
            .I2(n11280), .I3(rd_addr_r_c[2]), .O(n12959));
    defparam rd_addr_r_1__bdd_4_lut_11025.LUT_INIT = 16'he4aa;
    SB_LUT4 i3450_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_1_9 ), .O(n4833));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3450_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13619_bdd_4_lut (.I0(n13619), .I1(\REG.mem_25_8 ), .I2(\REG.mem_24_8 ), 
            .I3(rd_addr_r_c[1]), .O(n13622));
    defparam n13619_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4583_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_60_12 ), .O(n5966));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4583_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4582_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_60_11 ), .O(n5965));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4582_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4581_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_60_10 ), .O(n5964));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4581_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3484_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_1_14 ), .O(n4867));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3484_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3522_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_1_7 ), .O(n4905));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3522_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12959_bdd_4_lut (.I0(n12959), .I1(n11253), .I2(n11252), .I3(rd_addr_r_c[2]), 
            .O(n12962));
    defparam n12959_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3531_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_1_6 ), .O(n4914));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3531_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4087_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_33_12 ), .O(n5470));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4087_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1310_1311 (.Q(\REG.mem_13_8 ), .C(FIFO_CLK_c), .D(n5130));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4580_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_60_9 ), .O(n5963));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4580_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4579_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_60_8 ), .O(n5962));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4579_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3449_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_1_15 ), .O(n4832));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3449_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11555 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_0 ), 
            .I2(\REG.mem_55_0 ), .I3(rd_addr_r_c[1]), .O(n13613));
    defparam rd_addr_r_0__bdd_4_lut_11555.LUT_INIT = 16'he4aa;
    SB_LUT4 i4578_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_60_7 ), .O(n5961));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4578_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13613_bdd_4_lut (.I0(n13613), .I1(\REG.mem_53_0 ), .I2(\REG.mem_52_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11977));
    defparam n13613_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4577_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_60_6 ), .O(n5960));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4577_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1307_1308 (.Q(\REG.mem_13_7 ), .C(FIFO_CLK_c), .D(n5129));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1304_1305 (.Q(\REG.mem_13_6 ), .C(FIFO_CLK_c), .D(n5128));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1301_1302 (.Q(\REG.mem_13_5 ), .C(FIFO_CLK_c), .D(n5127));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1298_1299 (.Q(\REG.mem_13_4 ), .C(FIFO_CLK_c), .D(n5126));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4576_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_60_5 ), .O(n5959));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4576_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4575_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_60_4 ), .O(n5958));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4575_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1295_1296 (.Q(\REG.mem_13_3 ), .C(FIFO_CLK_c), .D(n5125));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11005 (.I0(rd_addr_r_c[1]), .I1(n11210), 
            .I2(n11211), .I3(rd_addr_r_c[2]), .O(n12953));
    defparam rd_addr_r_1__bdd_4_lut_11005.LUT_INIT = 16'he4aa;
    SB_LUT4 i4574_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_60_3 ), .O(n5957));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4574_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12953_bdd_4_lut (.I0(n12953), .I1(n11187), .I2(n11186), .I3(rd_addr_r_c[2]), 
            .O(n12956));
    defparam n12953_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1292_1293 (.Q(\REG.mem_13_2 ), .C(FIFO_CLK_c), .D(n5124));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11650 (.I0(rd_addr_r_c[2]), .I1(n13298), 
            .I2(n12482), .I3(rd_addr_r_c[3]), .O(n13607));
    defparam rd_addr_r_2__bdd_4_lut_11650.LUT_INIT = 16'he4aa;
    SB_LUT4 n13607_bdd_4_lut (.I0(n13607), .I1(n11977), .I2(n11968), .I3(rd_addr_r_c[3]), 
            .O(n11983));
    defparam n13607_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1289_1290 (.Q(\REG.mem_13_1 ), .C(FIFO_CLK_c), .D(n5123));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3452_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_1_5 ), .O(n4835));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3452_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3454_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_1_4 ), .O(n4837));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3454_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11550 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_8 ), 
            .I2(\REG.mem_11_8 ), .I3(rd_addr_r_c[1]), .O(n13601));
    defparam rd_addr_r_0__bdd_4_lut_11550.LUT_INIT = 16'he4aa;
    SB_LUT4 i10033_3_lut (.I0(\REG.mem_22_14 ), .I1(\REG.mem_23_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11871));
    defparam i10033_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1286_1287 (.Q(\REG.mem_13_0 ), .C(FIFO_CLK_c), .D(n5122));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1235_1236 (.Q(\REG.mem_12_15 ), .C(FIFO_CLK_c), .D(n5121));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1232_1233 (.Q(\REG.mem_12_14 ), .C(FIFO_CLK_c), .D(n5120));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4573_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_60_2 ), .O(n5956));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4573_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1229_1230 (.Q(\REG.mem_12_13 ), .C(FIFO_CLK_c), .D(n5119));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1226_1227 (.Q(\REG.mem_12_12 ), .C(FIFO_CLK_c), .D(n5118));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3478_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_1_3 ), .O(n4861));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3478_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10524 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_6 ), 
            .I2(\REG.mem_35_6 ), .I3(rd_addr_r_c[1]), .O(n12371));
    defparam rd_addr_r_0__bdd_4_lut_10524.LUT_INIT = 16'he4aa;
    SB_LUT4 i3485_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_1_2 ), .O(n4868));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3485_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11010 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_9 ), 
            .I2(\REG.mem_3_9 ), .I3(rd_addr_r_c[1]), .O(n12947));
    defparam rd_addr_r_0__bdd_4_lut_11010.LUT_INIT = 16'he4aa;
    SB_LUT4 n13601_bdd_4_lut (.I0(n13601), .I1(\REG.mem_9_8 ), .I2(\REG.mem_8_8 ), 
            .I3(rd_addr_r_c[1]), .O(n13604));
    defparam n13601_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1223_1224 (.Q(\REG.mem_12_11 ), .C(FIFO_CLK_c), .D(n5117));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12947_bdd_4_lut (.I0(n12947), .I1(\REG.mem_1_9 ), .I2(\REG.mem_0_9 ), 
            .I3(rd_addr_r_c[1]), .O(n11122));
    defparam n12947_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9162_3_lut (.I0(\REG.mem_8_6 ), .I1(\REG.mem_9_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11000));
    defparam i9162_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1220_1221 (.Q(\REG.mem_12_10 ), .C(FIFO_CLK_c), .D(n5116));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9163_3_lut (.I0(\REG.mem_10_6 ), .I1(\REG.mem_11_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11001));
    defparam i9163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4572_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_60_1 ), .O(n5955));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4572_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11115 (.I0(rd_addr_r_c[2]), .I1(n11272), 
            .I2(n12452), .I3(rd_addr_r_c[3]), .O(n12941));
    defparam rd_addr_r_2__bdd_4_lut_11115.LUT_INIT = 16'he4aa;
    SB_LUT4 i3496_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_1_1 ), .O(n4879));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3496_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4571_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_60_0 ), .O(n5954));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4571_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10032_3_lut (.I0(\REG.mem_20_14 ), .I1(\REG.mem_21_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11870));
    defparam i10032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12941_bdd_4_lut (.I0(n12941), .I1(n11197), .I2(n11110), .I3(rd_addr_r_c[3]), 
            .O(n11704));
    defparam n12941_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3501_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_1_0 ), .O(n4884));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3501_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12287_bdd_4_lut (.I0(n12287), .I1(n11419), .I2(n11389), .I3(rd_addr_r_c[3]), 
            .O(n12290));
    defparam n12287_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i61_2_lut_3_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n61_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i61_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i94_2_lut_3_lut_4_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n53));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i94_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i93_2_lut_3_lut_4_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n21));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i93_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11565 (.I0(rd_addr_r_c[1]), .I1(n11432), 
            .I2(n11433), .I3(rd_addr_r_c[2]), .O(n13595));
    defparam rd_addr_r_1__bdd_4_lut_11565.LUT_INIT = 16'he4aa;
    SB_LUT4 n12371_bdd_4_lut (.I0(n12371), .I1(\REG.mem_33_6 ), .I2(\REG.mem_32_6 ), 
            .I3(rd_addr_r_c[1]), .O(n12374));
    defparam n12371_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i13_2_lut_3_lut_4_lut (.I0(wr_sig_mv_w), .I1(wr_addr_r[0]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[1]), .O(n13));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i13_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i3517_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_1_8 ), .O(n4900));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3517_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10995 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_1 ), 
            .I2(\REG.mem_59_1 ), .I3(rd_addr_r_c[1]), .O(n12935));
    defparam rd_addr_r_0__bdd_4_lut_10995.LUT_INIT = 16'he4aa;
    SB_DFF i1217_1218 (.Q(\REG.mem_12_9 ), .C(FIFO_CLK_c), .D(n5115));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1214_1215 (.Q(\REG.mem_12_8 ), .C(FIFO_CLK_c), .D(n5114));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1211_1212 (.Q(\REG.mem_12_7 ), .C(FIFO_CLK_c), .D(n5113));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i14_2_lut_3_lut_4_lut (.I0(wr_sig_mv_w), .I1(wr_addr_r[0]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[1]), .O(n14));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i14_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 n12935_bdd_4_lut (.I0(n12935), .I1(\REG.mem_57_1 ), .I2(\REG.mem_56_1 ), 
            .I3(rd_addr_r_c[1]), .O(n12938));
    defparam n12935_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4561_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_59_15 ), .O(n5944));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4561_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13595_bdd_4_lut (.I0(n13595), .I1(n11421), .I2(n11420), .I3(rd_addr_r_c[2]), 
            .O(n11514));
    defparam n13595_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4560_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_59_14 ), .O(n5943));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4560_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i2_2_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_w[2]), 
            .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[1] ), .O(wr_grey_w[1]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i2_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11545 (.I0(rd_addr_r_c[2]), .I1(n11440), 
            .I2(n11482), .I3(rd_addr_r_c[3]), .O(n13589));
    defparam rd_addr_r_2__bdd_4_lut_11545.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i3_2_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_w[2]), 
            .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[3] ), .O(wr_grey_w[2]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i3_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_DFF i1208_1209 (.Q(\REG.mem_12_6 ), .C(FIFO_CLK_c), .D(n5112));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4661_2_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_w[2]), 
            .I2(wr_sig_mv_w), .I3(reset_per_frame), .O(n6044));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i4661_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 i4559_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_59_13 ), .O(n5942));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4559_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4086_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_33_11 ), .O(n5469));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4086_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4558_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_59_12 ), .O(n5941));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4558_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4557_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_59_11 ), .O(n5940));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4557_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4556_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_59_10 ), .O(n5939));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4556_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13589_bdd_4_lut (.I0(n13589), .I1(n12398), .I2(n13184), .I3(rd_addr_r_c[3]), 
            .O(n11989));
    defparam n13589_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i100_2_lut_3_lut (.I0(n35), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n50));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i100_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10985 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_11 ), 
            .I2(\REG.mem_51_11 ), .I3(rd_addr_r_c[1]), .O(n12929));
    defparam rd_addr_r_0__bdd_4_lut_10985.LUT_INIT = 16'he4aa;
    SB_DFF i1205_1206 (.Q(\REG.mem_12_5 ), .C(FIFO_CLK_c), .D(n5111));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4555_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_59_9 ), .O(n5938));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4555_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4554_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_59_8 ), .O(n5937));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4554_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i99_2_lut_3_lut (.I0(n35), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n18));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i99_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i9718_3_lut (.I0(\REG.mem_6_12 ), .I1(\REG.mem_7_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11556));
    defparam i9718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4553_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_59_7 ), .O(n5936));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4553_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1202_1203 (.Q(\REG.mem_12_4 ), .C(FIFO_CLK_c), .D(n5110));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1199_1200 (.Q(\REG.mem_12_3 ), .C(FIFO_CLK_c), .D(n5109));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4552_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_59_6 ), .O(n5935));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4552_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4551_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_59_5 ), .O(n5934));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4551_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4550_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_59_4 ), .O(n5933));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4550_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4549_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_59_3 ), .O(n5932));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4549_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1196_1197 (.Q(\REG.mem_12_2 ), .C(FIFO_CLK_c), .D(n5108));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i4_2_lut_4_lut (.I0(wr_addr_r[4]), .I1(wr_addr_p1_w[4]), 
            .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[3] ), .O(wr_grey_w[3]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i4_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 n12929_bdd_4_lut (.I0(n12929), .I1(\REG.mem_49_11 ), .I2(\REG.mem_48_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11710));
    defparam n12929_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9717_3_lut (.I0(\REG.mem_4_12 ), .I1(\REG.mem_5_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11555));
    defparam i9717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4548_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_59_2 ), .O(n5931));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4548_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10519 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_2 ), 
            .I2(\REG.mem_11_2 ), .I3(rd_addr_r_c[1]), .O(n12365));
    defparam rd_addr_r_0__bdd_4_lut_10519.LUT_INIT = 16'he4aa;
    SB_LUT4 i4547_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_59_1 ), .O(n5930));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4547_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i5_2_lut_4_lut (.I0(wr_addr_r[4]), .I1(wr_addr_p1_w[4]), 
            .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[5] ), .O(wr_grey_w[4]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i5_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4546_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_59_0 ), .O(n5929));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4546_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1193_1194 (.Q(\REG.mem_12_1 ), .C(FIFO_CLK_c), .D(n5107));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12365_bdd_4_lut (.I0(n12365), .I1(\REG.mem_9_2 ), .I2(\REG.mem_8_2 ), 
            .I3(rd_addr_r_c[1]), .O(n12368));
    defparam n12365_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i92_2_lut_3_lut_4_lut (.I0(n20_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n54));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i92_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i91_2_lut_3_lut_4_lut (.I0(n20_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n22));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i91_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i4659_2_lut_4_lut (.I0(wr_addr_r[4]), .I1(wr_addr_p1_w[4]), 
            .I2(wr_sig_mv_w), .I3(reset_per_frame), .O(n6042));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i4659_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 i4085_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_33_10 ), .O(n5468));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4085_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10980 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_0 ), 
            .I2(\REG.mem_15_0 ), .I3(rd_addr_r_c[1]), .O(n12923));
    defparam rd_addr_r_0__bdd_4_lut_10980.LUT_INIT = 16'he4aa;
    SB_DFF i1190_1191 (.Q(\REG.mem_12_0 ), .C(FIFO_CLK_c), .D(n5106));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i4_2_lut_4_lut (.I0(rd_addr_r_c[4]), 
            .I1(rd_addr_p1_w[4]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_498[3] ), 
            .O(rd_grey_w[3]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i4_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 n12923_bdd_4_lut (.I0(n12923), .I1(\REG.mem_13_0 ), .I2(\REG.mem_12_0 ), 
            .I3(rd_addr_r_c[1]), .O(n12926));
    defparam n12923_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9256_3_lut (.I0(\REG.mem_14_6 ), .I1(\REG.mem_15_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11094));
    defparam i9256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11660 (.I0(rd_addr_r_c[3]), .I1(n13022), 
            .I2(n11514), .I3(rd_addr_r_c[4]), .O(n13583));
    defparam rd_addr_r_3__bdd_4_lut_11660.LUT_INIT = 16'he4aa;
    SB_LUT4 i9255_3_lut (.I0(\REG.mem_12_6 ), .I1(\REG.mem_13_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11093));
    defparam i9255_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1139_1140 (.Q(\REG.mem_11_15 ), .C(FIFO_CLK_c), .D(n5105));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1136_1137 (.Q(\REG.mem_11_14 ), .C(FIFO_CLK_c), .D(n5104));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1133_1134 (.Q(\REG.mem_11_13 ), .C(FIFO_CLK_c), .D(n5103));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1130_1131 (.Q(\REG.mem_11_12 ), .C(FIFO_CLK_c), .D(n5102));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1127_1128 (.Q(\REG.mem_11_11 ), .C(FIFO_CLK_c), .D(n5101));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1124_1125 (.Q(\REG.mem_11_10 ), .C(FIFO_CLK_c), .D(n5100));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1121_1122 (.Q(\REG.mem_11_9 ), .C(FIFO_CLK_c), .D(n5099));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1118_1119 (.Q(\REG.mem_11_8 ), .C(FIFO_CLK_c), .D(n5098));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i140_141 (.Q(\REG.mem_1_2 ), .C(FIFO_CLK_c), .D(n4868));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i176_177 (.Q(\REG.mem_1_14 ), .C(FIFO_CLK_c), .D(n4867));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wr_addr_r__i0 (.Q(wr_addr_r[0]), .C(FIFO_CLK_c), .D(n4866));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF i143_144 (.Q(\REG.mem_1_3 ), .C(FIFO_CLK_c), .D(n4861));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10975 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_12 ), 
            .I2(\REG.mem_43_12 ), .I3(rd_addr_r_c[1]), .O(n12917));
    defparam rd_addr_r_0__bdd_4_lut_10975.LUT_INIT = 16'he4aa;
    SB_LUT4 n13583_bdd_4_lut (.I0(n13583), .I1(n11493), .I2(n11492), .I3(rd_addr_r_c[4]), 
            .O(n13586));
    defparam n13583_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1115_1116 (.Q(\REG.mem_11_7 ), .C(FIFO_CLK_c), .D(n5097));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11540 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_6 ), 
            .I2(\REG.mem_23_6 ), .I3(rd_addr_r_c[1]), .O(n13577));
    defparam rd_addr_r_0__bdd_4_lut_11540.LUT_INIT = 16'he4aa;
    SB_DFF i1112_1113 (.Q(\REG.mem_11_6 ), .C(FIFO_CLK_c), .D(n5096));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1109_1110 (.Q(\REG.mem_11_5 ), .C(FIFO_CLK_c), .D(n5095));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1106_1107 (.Q(\REG.mem_11_4 ), .C(FIFO_CLK_c), .D(n5094));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1103_1104 (.Q(\REG.mem_11_3 ), .C(FIFO_CLK_c), .D(n5093));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1100_1101 (.Q(\REG.mem_11_2 ), .C(FIFO_CLK_c), .D(n5092));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1097_1098 (.Q(\REG.mem_11_1 ), .C(FIFO_CLK_c), .D(n5091));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1094_1095 (.Q(\REG.mem_11_0 ), .C(FIFO_CLK_c), .D(n5090));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1043_1044 (.Q(\REG.mem_10_15 ), .C(FIFO_CLK_c), .D(n5089));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12917_bdd_4_lut (.I0(n12917), .I1(\REG.mem_41_12 ), .I2(\REG.mem_40_12 ), 
            .I3(rd_addr_r_c[1]), .O(n12920));
    defparam n12917_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1040_1041 (.Q(\REG.mem_10_14 ), .C(FIFO_CLK_c), .D(n5088));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10970 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_0 ), 
            .I2(\REG.mem_19_0 ), .I3(rd_addr_r_c[1]), .O(n12911));
    defparam rd_addr_r_0__bdd_4_lut_10970.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i5_2_lut_4_lut (.I0(rd_addr_r_c[4]), 
            .I1(rd_addr_p1_w[4]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_498[5] ), 
            .O(rd_grey_w[4]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i5_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 n13577_bdd_4_lut (.I0(n13577), .I1(\REG.mem_21_6 ), .I2(\REG.mem_20_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11197));
    defparam n13577_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12911_bdd_4_lut (.I0(n12911), .I1(\REG.mem_17_0 ), .I2(\REG.mem_16_0 ), 
            .I3(rd_addr_r_c[1]), .O(n12914));
    defparam n12911_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1037_1038 (.Q(\REG.mem_10_13 ), .C(FIFO_CLK_c), .D(n5087));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1034_1035 (.Q(\REG.mem_10_12 ), .C(FIFO_CLK_c), .D(n5086));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1031_1032 (.Q(\REG.mem_10_11 ), .C(FIFO_CLK_c), .D(n5085));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1028_1029 (.Q(\REG.mem_10_10 ), .C(FIFO_CLK_c), .D(n5084));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1025_1026 (.Q(\REG.mem_10_9 ), .C(FIFO_CLK_c), .D(n5083));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1022_1023 (.Q(\REG.mem_10_8 ), .C(FIFO_CLK_c), .D(n5082));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1019_1020 (.Q(\REG.mem_10_7 ), .C(FIFO_CLK_c), .D(n5081));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1016_1017 (.Q(\REG.mem_10_6 ), .C(FIFO_CLK_c), .D(n5080));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4539_2_lut_4_lut (.I0(rd_addr_r_c[4]), .I1(rd_addr_p1_w[4]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n5922));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4539_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 rd_addr_r_6__I_0_i6_3_lut (.I0(rd_addr_r_c[5]), .I1(rd_addr_p1_w[5]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_6__N_498[5] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_6__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1013_1014 (.Q(\REG.mem_10_5 ), .C(FIFO_CLK_c), .D(n5079));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10965 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_1 ), 
            .I2(\REG.mem_11_1 ), .I3(rd_addr_r_c[1]), .O(n12905));
    defparam rd_addr_r_0__bdd_4_lut_10965.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i6_2_lut_4_lut (.I0(\rd_addr_r[6] ), 
            .I1(rd_addr_p1_w[6]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_498[5] ), 
            .O(rd_grey_w[5]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i6_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4537_2_lut_4_lut (.I0(\rd_addr_r[6] ), .I1(rd_addr_p1_w[6]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n5920));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4537_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11520 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_6 ), 
            .I2(\REG.mem_51_6 ), .I3(rd_addr_r_c[1]), .O(n13571));
    defparam rd_addr_r_0__bdd_4_lut_11520.LUT_INIT = 16'he4aa;
    SB_LUT4 i4536_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_58_15 ), .O(n5919));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4536_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12905_bdd_4_lut (.I0(n12905), .I1(\REG.mem_9_1 ), .I2(\REG.mem_8_1 ), 
            .I3(rd_addr_r_c[1]), .O(n11302));
    defparam n12905_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4084_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_33_9 ), .O(n5467));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4084_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13571_bdd_4_lut (.I0(n13571), .I1(\REG.mem_49_6 ), .I2(\REG.mem_48_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11530));
    defparam n13571_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4535_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_58_14 ), .O(n5918));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4535_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10960 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_11 ), 
            .I2(\REG.mem_55_11 ), .I3(rd_addr_r_c[1]), .O(n12899));
    defparam rd_addr_r_0__bdd_4_lut_10960.LUT_INIT = 16'he4aa;
    SB_LUT4 i4534_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_58_13 ), .O(n5917));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4534_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4533_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_58_12 ), .O(n5916));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4533_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4532_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_58_11 ), .O(n5915));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4532_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11530 (.I0(rd_addr_r_c[2]), .I1(n13226), 
            .I2(n12836), .I3(rd_addr_r_c[3]), .O(n13565));
    defparam rd_addr_r_2__bdd_4_lut_11530.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_6__I_0_i4_3_lut (.I0(rd_addr_r_c[3]), .I1(rd_addr_p1_w[3]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_6__N_498[3] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_6__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13565_bdd_4_lut (.I0(n13565), .I1(n13418), .I2(n11500), .I3(rd_addr_r_c[3]), 
            .O(n11995));
    defparam n13565_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4531_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_58_10 ), .O(n5914));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4531_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_6__I_0_i3_3_lut (.I0(rd_addr_r_c[2]), .I1(rd_addr_p1_w[2]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_6__N_498[2] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_6__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4530_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_58_9 ), .O(n5913));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4530_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4529_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_58_8 ), .O(n5912));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4529_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4528_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_58_7 ), .O(n5911));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4528_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12899_bdd_4_lut (.I0(n12899), .I1(\REG.mem_53_11 ), .I2(\REG.mem_52_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11719));
    defparam n12899_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i88_2_lut_3_lut (.I0(n23_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n56));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i88_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i4527_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_58_6 ), .O(n5910));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4527_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4526_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_58_5 ), .O(n5909));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4526_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i87_2_lut_3_lut (.I0(n23_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n24));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i87_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i4083_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_33_8 ), .O(n5466));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4083_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10955 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_3 ), 
            .I2(\REG.mem_59_3 ), .I3(rd_addr_r_c[1]), .O(n12893));
    defparam rd_addr_r_0__bdd_4_lut_10955.LUT_INIT = 16'he4aa;
    SB_LUT4 i4525_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_58_4 ), .O(n5908));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4525_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4524_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_58_3 ), .O(n5907));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4524_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4523_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_58_2 ), .O(n5906));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4523_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12893_bdd_4_lut (.I0(n12893), .I1(\REG.mem_57_3 ), .I2(\REG.mem_56_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11125));
    defparam n12893_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_11630 (.I0(rd_addr_r_c[4]), .I1(n12554), 
            .I2(n11983), .I3(rd_addr_r_c[5]), .O(n13559));
    defparam rd_addr_r_4__bdd_4_lut_11630.LUT_INIT = 16'he4aa;
    SB_LUT4 n13559_bdd_4_lut (.I0(n13559), .I1(n13094), .I2(n11575), .I3(rd_addr_r_c[5]), 
            .O(\REG.out_raw_31__N_559 [0]));
    defparam n13559_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4522_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_58_1 ), .O(n5905));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4522_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1010_1011 (.Q(\REG.mem_10_4 ), .C(FIFO_CLK_c), .D(n5078));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4521_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_58_0 ), .O(n5904));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4521_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11515 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_3 ), 
            .I2(\REG.mem_15_3 ), .I3(rd_addr_r_c[1]), .O(n13553));
    defparam rd_addr_r_0__bdd_4_lut_11515.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i90_2_lut_3_lut_4_lut (.I0(n18_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n55));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i90_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i89_2_lut_3_lut_4_lut (.I0(n18_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n23));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i89_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_DFF i1007_1008 (.Q(\REG.mem_10_3 ), .C(FIFO_CLK_c), .D(n5077));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i120_2_lut_3_lut (.I0(n23_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n40));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i120_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i119_2_lut_3_lut (.I0(n23_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n8));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i119_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10950 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_5 ), 
            .I2(\REG.mem_35_5 ), .I3(rd_addr_r_c[1]), .O(n12887));
    defparam rd_addr_r_0__bdd_4_lut_10950.LUT_INIT = 16'he4aa;
    SB_LUT4 n13553_bdd_4_lut (.I0(n13553), .I1(\REG.mem_13_3 ), .I2(\REG.mem_12_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11056));
    defparam n13553_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12887_bdd_4_lut (.I0(n12887), .I1(\REG.mem_33_5 ), .I2(\REG.mem_32_5 ), 
            .I3(rd_addr_r_c[1]), .O(n12890));
    defparam n12887_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i23_2_lut_3_lut (.I0(n12_adj_33), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n23_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i23_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_11505 (.I0(rd_addr_r_c[4]), .I1(n11989), 
            .I2(n11995), .I3(rd_addr_r_c[5]), .O(n13547));
    defparam rd_addr_r_4__bdd_4_lut_11505.LUT_INIT = 16'he4aa;
    SB_DFF i1004_1005 (.Q(\REG.mem_10_2 ), .C(FIFO_CLK_c), .D(n5076));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1001_1002 (.Q(\REG.mem_10_1 ), .C(FIFO_CLK_c), .D(n5075));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10514 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_7 ), 
            .I2(\REG.mem_23_7 ), .I3(rd_addr_r_c[1]), .O(n12359));
    defparam rd_addr_r_0__bdd_4_lut_10514.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i40_2_lut_3_lut_4_lut (.I0(n12_adj_33), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n40_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i40_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 n13547_bdd_4_lut (.I0(n13547), .I1(n11914), .I2(n12314), .I3(rd_addr_r_c[5]), 
            .O(\REG.out_raw_31__N_559 [13]));
    defparam n13547_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i39_2_lut_3_lut_4_lut (.I0(n12_adj_33), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n39));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i39_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11060 (.I0(rd_addr_r_c[3]), .I1(n12866), 
            .I2(n11256), .I3(rd_addr_r_c[4]), .O(n12881));
    defparam rd_addr_r_3__bdd_4_lut_11060.LUT_INIT = 16'he4aa;
    SB_LUT4 n12881_bdd_4_lut (.I0(n12881), .I1(n11250), .I2(n11249), .I3(rd_addr_r_c[4]), 
            .O(n12884));
    defparam n12881_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i998_999 (.Q(\REG.mem_10_0 ), .C(FIFO_CLK_c), .D(n5074));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11500 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_6 ), 
            .I2(\REG.mem_55_6 ), .I3(rd_addr_r_c[1]), .O(n13541));
    defparam rd_addr_r_0__bdd_4_lut_11500.LUT_INIT = 16'he4aa;
    SB_LUT4 n13541_bdd_4_lut (.I0(n13541), .I1(\REG.mem_53_6 ), .I2(\REG.mem_52_6 ), 
            .I3(rd_addr_r_c[1]), .O(n11545));
    defparam n13541_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11000 (.I0(rd_addr_r_c[1]), .I1(n11234), 
            .I2(n11235), .I3(rd_addr_r_c[2]), .O(n12875));
    defparam rd_addr_r_1__bdd_4_lut_11000.LUT_INIT = 16'he4aa;
    SB_DFF i947_948 (.Q(\REG.mem_9_15 ), .C(FIFO_CLK_c), .D(n5073));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4082_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_33_7 ), .O(n5465));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4082_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4501_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_56_15 ), .O(n5884));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4501_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4500_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_56_14 ), .O(n5883));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4500_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4499_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_56_13 ), .O(n5882));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4499_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4498_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_56_12 ), .O(n5881));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4498_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11490 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_3 ), 
            .I2(\REG.mem_19_3 ), .I3(rd_addr_r_c[1]), .O(n13535));
    defparam rd_addr_r_0__bdd_4_lut_11490.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10484 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_7 ), 
            .I2(\REG.mem_27_7 ), .I3(rd_addr_r_c[1]), .O(n12323));
    defparam rd_addr_r_0__bdd_4_lut_10484.LUT_INIT = 16'he4aa;
    SB_DFF i944_945 (.Q(\REG.mem_9_14 ), .C(FIFO_CLK_c), .D(n5072));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12875_bdd_4_lut (.I0(n12875), .I1(n11226), .I2(n11225), .I3(rd_addr_r_c[2]), 
            .O(n12878));
    defparam n12875_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4497_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_56_11 ), .O(n5880));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4497_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13535_bdd_4_lut (.I0(n13535), .I1(\REG.mem_17_3 ), .I2(\REG.mem_16_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11059));
    defparam n13535_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i20_2_lut (.I0(n11), .I1(wr_addr_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n20_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i20_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4496_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_56_10 ), .O(n5879));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4496_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i146_147 (.Q(\REG.mem_1_4 ), .C(FIFO_CLK_c), .D(n4837));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4495_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_56_9 ), .O(n5878));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4495_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10935 (.I0(rd_addr_r_c[1]), .I1(n11213), 
            .I2(n11214), .I3(rd_addr_r_c[2]), .O(n12869));
    defparam rd_addr_r_1__bdd_4_lut_10935.LUT_INIT = 16'he4aa;
    SB_LUT4 i4494_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_56_8 ), .O(n5877));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4494_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4493_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_56_7 ), .O(n5876));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4493_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4492_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_56_6 ), .O(n5875));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4492_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i941_942 (.Q(\REG.mem_9_13 ), .C(FIFO_CLK_c), .D(n5071));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11525 (.I0(rd_addr_r_c[3]), .I1(n12722), 
            .I2(n11052), .I3(rd_addr_r_c[4]), .O(n13529));
    defparam rd_addr_r_3__bdd_4_lut_11525.LUT_INIT = 16'he4aa;
    SB_DFF i938_939 (.Q(\REG.mem_9_12 ), .C(FIFO_CLK_c), .D(n5070));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4491_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_56_5 ), .O(n5874));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4491_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9672_3_lut (.I0(\REG.mem_56_7 ), .I1(\REG.mem_57_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11510));
    defparam i9672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12359_bdd_4_lut (.I0(n12359), .I1(\REG.mem_21_7 ), .I2(\REG.mem_20_7 ), 
            .I3(rd_addr_r_c[1]), .O(n12362));
    defparam n12359_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12869_bdd_4_lut (.I0(n12869), .I1(n11208), .I2(n11207), .I3(rd_addr_r_c[2]), 
            .O(n12872));
    defparam n12869_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9673_3_lut (.I0(\REG.mem_58_7 ), .I1(\REG.mem_59_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11511));
    defparam i9673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10930 (.I0(rd_addr_r_c[1]), .I1(n11189), 
            .I2(n11190), .I3(rd_addr_r_c[2]), .O(n12863));
    defparam rd_addr_r_1__bdd_4_lut_10930.LUT_INIT = 16'he4aa;
    SB_DFF i935_936 (.Q(\REG.mem_9_11 ), .C(FIFO_CLK_c), .D(n5069));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4490_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_56_4 ), .O(n5873));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4490_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12863_bdd_4_lut (.I0(n12863), .I1(n11178), .I2(n11177), .I3(rd_addr_r_c[2]), 
            .O(n12866));
    defparam n12863_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4489_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_56_3 ), .O(n5872));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4489_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4488_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_56_2 ), .O(n5871));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4488_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4487_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_56_1 ), .O(n5870));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4487_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_33 (.I0(DEBUG_3_c), .I1(get_next_word), .I2(GND_net), 
            .I3(GND_net), .O(rd_fifo_en_w));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i1_2_lut_adj_33.LUT_INIT = 16'h4444;
    SB_LUT4 n13529_bdd_4_lut (.I0(n13529), .I1(n11028), .I2(n11027), .I3(rd_addr_r_c[4]), 
            .O(n13532));
    defparam n13529_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4482_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_56_0 ), .O(n5865));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4482_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10509 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_15 ), 
            .I2(\REG.mem_47_15 ), .I3(rd_addr_r_c[1]), .O(n12353));
    defparam rd_addr_r_0__bdd_4_lut_10509.LUT_INIT = 16'he4aa;
    SB_DFF i149_150 (.Q(\REG.mem_1_5 ), .C(FIFO_CLK_c), .D(n4835));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i932_933 (.Q(\REG.mem_9_10 ), .C(FIFO_CLK_c), .D(n5068));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i929_930 (.Q(\REG.mem_9_9 ), .C(FIFO_CLK_c), .D(n5067));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10945 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_11 ), 
            .I2(\REG.mem_59_11 ), .I3(rd_addr_r_c[1]), .O(n12857));
    defparam rd_addr_r_0__bdd_4_lut_10945.LUT_INIT = 16'he4aa;
    SB_LUT4 n12857_bdd_4_lut (.I0(n12857), .I1(\REG.mem_57_11 ), .I2(\REG.mem_56_11 ), 
            .I3(rd_addr_r_c[1]), .O(n11722));
    defparam n12857_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i926_927 (.Q(\REG.mem_9_8 ), .C(FIFO_CLK_c), .D(n5066));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9694_3_lut (.I0(\REG.mem_62_7 ), .I1(\REG.mem_63_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11532));
    defparam i9694_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i923_924 (.Q(\REG.mem_9_7 ), .C(FIFO_CLK_c), .D(n5065));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11535 (.I0(rd_addr_r_c[1]), .I1(n11435), 
            .I2(n11436), .I3(rd_addr_r_c[2]), .O(n13523));
    defparam rd_addr_r_1__bdd_4_lut_11535.LUT_INIT = 16'he4aa;
    SB_LUT4 n13523_bdd_4_lut (.I0(n13523), .I1(n11427), .I2(n11426), .I3(rd_addr_r_c[2]), 
            .O(n11550));
    defparam n13523_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9693_3_lut (.I0(\REG.mem_60_7 ), .I1(\REG.mem_61_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11531));
    defparam i9693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i53_2_lut_3_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n53_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i53_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i86_2_lut_3_lut_4_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n57));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i86_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11485 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_3 ), 
            .I2(\REG.mem_23_3 ), .I3(rd_addr_r_c[1]), .O(n13517));
    defparam rd_addr_r_0__bdd_4_lut_11485.LUT_INIT = 16'he4aa;
    SB_DFF i920_921 (.Q(\REG.mem_9_6 ), .C(FIFO_CLK_c), .D(n5064));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13517_bdd_4_lut (.I0(n13517), .I1(\REG.mem_21_3 ), .I2(\REG.mem_20_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11065));
    defparam n13517_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i85_2_lut_3_lut_4_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n25));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i85_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i4081_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_33_6 ), .O(n5464));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4081_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11470 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_14 ), 
            .I2(\REG.mem_51_14 ), .I3(rd_addr_r_c[1]), .O(n13511));
    defparam rd_addr_r_0__bdd_4_lut_11470.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i2_2_lut_4_lut (.I0(rd_addr_r_c[1]), 
            .I1(rd_addr_p1_w[1]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_498[2] ), 
            .O(rd_grey_w[1]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i2_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 n13511_bdd_4_lut (.I0(n13511), .I1(\REG.mem_49_14 ), .I2(\REG.mem_48_14 ), 
            .I3(rd_addr_r_c[1]), .O(n12010));
    defparam n13511_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i917_918 (.Q(\REG.mem_9_5 ), .C(FIFO_CLK_c), .D(n5063));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10920 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_0 ), 
            .I2(\REG.mem_23_0 ), .I3(rd_addr_r_c[1]), .O(n12851));
    defparam rd_addr_r_0__bdd_4_lut_10920.LUT_INIT = 16'he4aa;
    SB_LUT4 n12851_bdd_4_lut (.I0(n12851), .I1(\REG.mem_21_0 ), .I2(\REG.mem_20_0 ), 
            .I3(rd_addr_r_c[1]), .O(n12854));
    defparam n12851_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11465 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_14 ), 
            .I2(\REG.mem_55_14 ), .I3(rd_addr_r_c[1]), .O(n13505));
    defparam rd_addr_r_0__bdd_4_lut_11465.LUT_INIT = 16'he4aa;
    SB_LUT4 i4542_2_lut_4_lut (.I0(rd_addr_r_c[1]), .I1(rd_addr_p1_w[1]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n5925));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4542_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 n13505_bdd_4_lut (.I0(n13505), .I1(\REG.mem_53_14 ), .I2(\REG.mem_52_14 ), 
            .I3(rd_addr_r_c[1]), .O(n12016));
    defparam n13505_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i914_915 (.Q(\REG.mem_9_4 ), .C(FIFO_CLK_c), .D(n5062));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4080_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_33_5 ), .O(n5463));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4080_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_34 (.I0(rp_sync2_r[5]), .I1(rp_sync2_r[4]), .I2(rp_sync2_r[6]), 
            .I3(GND_net), .O(rp_sync_w[4]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i2_3_lut_adj_34.LUT_INIT = 16'h6969;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i1_2_lut_4_lut (.I0(rd_addr_r_c[1]), 
            .I1(rd_addr_p1_w[1]), .I2(rd_fifo_en_w), .I3(rd_addr_nxt_c_6__N_498[0]), 
            .O(rd_grey_w[0]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i1_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i1_2_lut_adj_35 (.I0(rp_sync2_r[3]), .I1(rp_sync_w[4]), .I2(GND_net), 
            .I3(GND_net), .O(rp_sync_w[3]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_adj_35.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_36 (.I0(rp_sync2_r[1]), .I1(rp_sync_w[2]), .I2(GND_net), 
            .I3(GND_net), .O(rp_sync_w[1]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_adj_36.LUT_INIT = 16'h6666;
    SB_LUT4 i3483_2_lut_4_lut (.I0(wr_addr_r[0]), .I1(wr_addr_p1_w[0]), 
            .I2(wr_sig_mv_w), .I3(reset_per_frame), .O(n4866));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i3483_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 rp_sync2_r_6__I_0_136_i1_2_lut (.I0(rp_sync2_r[5]), .I1(rp_sync2_r[6]), 
            .I2(GND_net), .I3(GND_net), .O(rp_sync_w[5]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam rp_sync2_r_6__I_0_136_i1_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i1_2_lut_4_lut (.I0(wr_addr_r[0]), .I1(wr_addr_p1_w[0]), 
            .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[1] ), .O(wr_grey_w[0]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i1_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_DFF i911_912 (.Q(\REG.mem_9_3 ), .C(FIFO_CLK_c), .D(n5061));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3561_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_0_0 ), .O(n4944));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3561_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3541_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_0_15 ), .O(n4924));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3541_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3542_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_0_14 ), .O(n4925));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3542_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3543_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_0_13 ), .O(n4926));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3543_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3544_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_0_12 ), .O(n4927));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3544_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3545_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_0_11 ), .O(n4928));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3545_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i908_909 (.Q(\REG.mem_9_2 ), .C(FIFO_CLK_c), .D(n5060));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i905_906 (.Q(\REG.mem_9_1 ), .C(FIFO_CLK_c), .D(n5059));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i902_903 (.Q(\REG.mem_9_0 ), .C(FIFO_CLK_c), .D(n5057));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i851_852 (.Q(\REG.mem_8_15 ), .C(FIFO_CLK_c), .D(n5056));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i848_849 (.Q(\REG.mem_8_14 ), .C(FIFO_CLK_c), .D(n5055));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i845_846 (.Q(\REG.mem_8_13 ), .C(FIFO_CLK_c), .D(n5054));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i842_843 (.Q(\REG.mem_8_12 ), .C(FIFO_CLK_c), .D(n5053));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i839_840 (.Q(\REG.mem_8_11 ), .C(FIFO_CLK_c), .D(n5052));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i836_837 (.Q(\REG.mem_8_10 ), .C(FIFO_CLK_c), .D(n5051));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i833_834 (.Q(\REG.mem_8_9 ), .C(FIFO_CLK_c), .D(n5050));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i830_831 (.Q(\REG.mem_8_8 ), .C(FIFO_CLK_c), .D(n5049));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i827_828 (.Q(\REG.mem_8_7 ), .C(FIFO_CLK_c), .D(n5048));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i824_825 (.Q(\REG.mem_8_6 ), .C(FIFO_CLK_c), .D(n5047));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i821_822 (.Q(\REG.mem_8_5 ), .C(FIFO_CLK_c), .D(n5046));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i818_819 (.Q(\REG.mem_8_4 ), .C(FIFO_CLK_c), .D(n5045));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i815_816 (.Q(\REG.mem_8_3 ), .C(FIFO_CLK_c), .D(n5044));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i812_813 (.Q(\REG.mem_8_2 ), .C(FIFO_CLK_c), .D(n5043));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i809_810 (.Q(\REG.mem_8_1 ), .C(FIFO_CLK_c), .D(n5042));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i806_807 (.Q(\REG.mem_8_0 ), .C(FIFO_CLK_c), .D(n5041));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i755_756 (.Q(\REG.mem_7_15 ), .C(FIFO_CLK_c), .D(n5040));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i752_753 (.Q(\REG.mem_7_14 ), .C(FIFO_CLK_c), .D(n5039));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i749_750 (.Q(\REG.mem_7_13 ), .C(FIFO_CLK_c), .D(n5038));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i746_747 (.Q(\REG.mem_7_12 ), .C(FIFO_CLK_c), .D(n5037));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i743_744 (.Q(\REG.mem_7_11 ), .C(FIFO_CLK_c), .D(n5036));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i740_741 (.Q(\REG.mem_7_10 ), .C(FIFO_CLK_c), .D(n5035));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i737_738 (.Q(\REG.mem_7_9 ), .C(FIFO_CLK_c), .D(n5034));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i734_735 (.Q(\REG.mem_7_8 ), .C(FIFO_CLK_c), .D(n5033));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i731_732 (.Q(\REG.mem_7_7 ), .C(FIFO_CLK_c), .D(n5032));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i728_729 (.Q(\REG.mem_7_6 ), .C(FIFO_CLK_c), .D(n5031));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i725_726 (.Q(\REG.mem_7_5 ), .C(FIFO_CLK_c), .D(n5030));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i722_723 (.Q(\REG.mem_7_4 ), .C(FIFO_CLK_c), .D(n5029));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i719_720 (.Q(\REG.mem_7_3 ), .C(FIFO_CLK_c), .D(n5028));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i716_717 (.Q(\REG.mem_7_2 ), .C(FIFO_CLK_c), .D(n5027));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i713_714 (.Q(\REG.mem_7_1 ), .C(FIFO_CLK_c), .D(n5026));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i710_711 (.Q(\REG.mem_7_0 ), .C(FIFO_CLK_c), .D(n5025));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i659_660 (.Q(\REG.mem_6_15 ), .C(FIFO_CLK_c), .D(n5024));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i656_657 (.Q(\REG.mem_6_14 ), .C(FIFO_CLK_c), .D(n5023));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i653_654 (.Q(\REG.mem_6_13 ), .C(FIFO_CLK_c), .D(n5022));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i650_651 (.Q(\REG.mem_6_12 ), .C(FIFO_CLK_c), .D(n5021));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i647_648 (.Q(\REG.mem_6_11 ), .C(FIFO_CLK_c), .D(n5020));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i644_645 (.Q(\REG.mem_6_10 ), .C(FIFO_CLK_c), .D(n5019));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i641_642 (.Q(\REG.mem_6_9 ), .C(FIFO_CLK_c), .D(n5018));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i638_639 (.Q(\REG.mem_6_8 ), .C(FIFO_CLK_c), .D(n5017));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i635_636 (.Q(\REG.mem_6_7 ), .C(FIFO_CLK_c), .D(n5016));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i632_633 (.Q(\REG.mem_6_6 ), .C(FIFO_CLK_c), .D(n5015));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i629_630 (.Q(\REG.mem_6_5 ), .C(FIFO_CLK_c), .D(n5014));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i626_627 (.Q(\REG.mem_6_4 ), .C(FIFO_CLK_c), .D(n5013));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i623_624 (.Q(\REG.mem_6_3 ), .C(FIFO_CLK_c), .D(n5012));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i620_621 (.Q(\REG.mem_6_2 ), .C(FIFO_CLK_c), .D(n5011));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i617_618 (.Q(\REG.mem_6_1 ), .C(FIFO_CLK_c), .D(n5010));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i614_615 (.Q(\REG.mem_6_0 ), .C(FIFO_CLK_c), .D(n5009));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i563_564 (.Q(\REG.mem_5_15 ), .C(FIFO_CLK_c), .D(n5008));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i560_561 (.Q(\REG.mem_5_14 ), .C(FIFO_CLK_c), .D(n5007));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i557_558 (.Q(\REG.mem_5_13 ), .C(FIFO_CLK_c), .D(n5006));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i554_555 (.Q(\REG.mem_5_12 ), .C(FIFO_CLK_c), .D(n5005));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i551_552 (.Q(\REG.mem_5_11 ), .C(FIFO_CLK_c), .D(n5004));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i548_549 (.Q(\REG.mem_5_10 ), .C(FIFO_CLK_c), .D(n5003));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i545_546 (.Q(\REG.mem_5_9 ), .C(FIFO_CLK_c), .D(n5002));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i542_543 (.Q(\REG.mem_5_8 ), .C(FIFO_CLK_c), .D(n5001));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i539_540 (.Q(\REG.mem_5_7 ), .C(FIFO_CLK_c), .D(n5000));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i536_537 (.Q(\REG.mem_5_6 ), .C(FIFO_CLK_c), .D(n4999));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i533_534 (.Q(\REG.mem_5_5 ), .C(FIFO_CLK_c), .D(n4998));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i530_531 (.Q(\REG.mem_5_4 ), .C(FIFO_CLK_c), .D(n4997));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i527_528 (.Q(\REG.mem_5_3 ), .C(FIFO_CLK_c), .D(n4996));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i524_525 (.Q(\REG.mem_5_2 ), .C(FIFO_CLK_c), .D(n4995));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i521_522 (.Q(\REG.mem_5_1 ), .C(FIFO_CLK_c), .D(n4994));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i518_519 (.Q(\REG.mem_5_0 ), .C(FIFO_CLK_c), .D(n4993));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i467_468 (.Q(\REG.mem_4_15 ), .C(FIFO_CLK_c), .D(n4992));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i464_465 (.Q(\REG.mem_4_14 ), .C(FIFO_CLK_c), .D(n4991));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i461_462 (.Q(\REG.mem_4_13 ), .C(FIFO_CLK_c), .D(n4990));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i458_459 (.Q(\REG.mem_4_12 ), .C(FIFO_CLK_c), .D(n4989));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i455_456 (.Q(\REG.mem_4_11 ), .C(FIFO_CLK_c), .D(n4988));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i452_453 (.Q(\REG.mem_4_10 ), .C(FIFO_CLK_c), .D(n4987));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i449_450 (.Q(\REG.mem_4_9 ), .C(FIFO_CLK_c), .D(n4986));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i446_447 (.Q(\REG.mem_4_8 ), .C(FIFO_CLK_c), .D(n4985));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i443_444 (.Q(\REG.mem_4_7 ), .C(FIFO_CLK_c), .D(n4984));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i440_441 (.Q(\REG.mem_4_6 ), .C(FIFO_CLK_c), .D(n4983));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i437_438 (.Q(\REG.mem_4_5 ), .C(FIFO_CLK_c), .D(n4982));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i434_435 (.Q(\REG.mem_4_4 ), .C(FIFO_CLK_c), .D(n4981));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i431_432 (.Q(\REG.mem_4_3 ), .C(FIFO_CLK_c), .D(n4980));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i428_429 (.Q(\REG.mem_4_2 ), .C(FIFO_CLK_c), .D(n4979));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i425_426 (.Q(\REG.mem_4_1 ), .C(FIFO_CLK_c), .D(n4978));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i422_423 (.Q(\REG.mem_4_0 ), .C(FIFO_CLK_c), .D(n4977));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i371_372 (.Q(\REG.mem_3_15 ), .C(FIFO_CLK_c), .D(n4976));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i368_369 (.Q(\REG.mem_3_14 ), .C(FIFO_CLK_c), .D(n4975));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i365_366 (.Q(\REG.mem_3_13 ), .C(FIFO_CLK_c), .D(n4974));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i362_363 (.Q(\REG.mem_3_12 ), .C(FIFO_CLK_c), .D(n4973));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i359_360 (.Q(\REG.mem_3_11 ), .C(FIFO_CLK_c), .D(n4972));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i356_357 (.Q(\REG.mem_3_10 ), .C(FIFO_CLK_c), .D(n4971));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i353_354 (.Q(\REG.mem_3_9 ), .C(FIFO_CLK_c), .D(n4970));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i350_351 (.Q(\REG.mem_3_8 ), .C(FIFO_CLK_c), .D(n4969));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12317_bdd_4_lut (.I0(n12317), .I1(n11143), .I2(n11122), .I3(rd_addr_r_c[3]), 
            .O(n12320));
    defparam n12317_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12353_bdd_4_lut (.I0(n12353), .I1(\REG.mem_45_15 ), .I2(\REG.mem_44_15 ), 
            .I3(rd_addr_r_c[1]), .O(n12356));
    defparam n12353_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3546_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_0_10 ), .O(n4929));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3546_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3547_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_0_9 ), .O(n4930));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3547_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11475 (.I0(rd_addr_r_c[1]), .I1(n11468), 
            .I2(n11469), .I3(rd_addr_r_c[2]), .O(n13499));
    defparam rd_addr_r_1__bdd_4_lut_11475.LUT_INIT = 16'he4aa;
    SB_LUT4 i9009_4_lut (.I0(wr_addr_r[1]), .I1(wr_addr_r[3]), .I2(rp_sync_w[1]), 
            .I3(rp_sync_w[3]), .O(n10845));
    defparam i9009_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 n13499_bdd_4_lut (.I0(n13499), .I1(n11457), .I2(n11456), .I3(rd_addr_r_c[2]), 
            .O(n11559));
    defparam n13499_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_p1_w_6__I_0_2_lut (.I0(wr_addr_p1_w[6]), .I1(rp_sync2_r[6]), 
            .I2(GND_net), .I3(GND_net), .O(full_max_w));   // src/fifo_dc_32_lut_gen.v(296[27:88])
    defparam wr_addr_p1_w_6__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10915 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_3 ), 
            .I2(\REG.mem_63_3 ), .I3(rd_addr_r_c[1]), .O(n12845));
    defparam rd_addr_r_0__bdd_4_lut_10915.LUT_INIT = 16'he4aa;
    SB_LUT4 i9013_4_lut (.I0(wr_addr_p1_w[4]), .I1(wr_addr_p1_w[1]), .I2(rp_sync_w[4]), 
            .I3(rp_sync_w[1]), .O(n10849));
    defparam i9013_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 i9045_4_lut (.I0(wr_addr_p1_w[5]), .I1(wr_addr_p1_w[3]), .I2(rp_sync_w[5]), 
            .I3(rp_sync_w[3]), .O(n10881));
    defparam i9045_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 i5_4_lut_adj_37 (.I0(wr_addr_p1_w[0]), .I1(n10849), .I2(full_max_w), 
            .I3(rp_sync_w[0]), .O(n12_adj_35));
    defparam i5_4_lut_adj_37.LUT_INIT = 16'h1020;
    SB_LUT4 wr_addr_r_5__I_0_i3_2_lut (.I0(wr_addr_r[2]), .I1(rp_sync_w[2]), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_36));   // src/fifo_dc_32_lut_gen.v(295[31:67])
    defparam wr_addr_r_5__I_0_i3_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i9110_4_lut (.I0(wr_addr_r[0]), .I1(n10845), .I2(n6_adj_37), 
            .I3(rp_sync_w[0]), .O(n10947));
    defparam i9110_4_lut.LUT_INIT = 16'hfefd;
    SB_LUT4 i10355_4_lut (.I0(wr_addr_p1_w[2]), .I1(n12_adj_35), .I2(n10881), 
            .I3(rp_sync_w[2]), .O(n12032));   // src/fifo_dc_32_lut_gen.v(300[45:114])
    defparam i10355_4_lut.LUT_INIT = 16'h0408;
    SB_LUT4 i10354_4_lut (.I0(wr_addr_r[4]), .I1(full_o), .I2(rp_sync_w[4]), 
            .I3(n3_adj_36), .O(n12033));   // src/fifo_dc_32_lut_gen.v(300[45:114])
    defparam i10354_4_lut.LUT_INIT = 16'h0048;
    SB_LUT4 full_nxt_c_I_6_4_lut (.I0(n12033), .I1(n12032), .I2(wr_sig_mv_w), 
            .I3(n10947), .O(full_nxt_c_N_626));   // src/fifo_dc_32_lut_gen.v(300[45:114])
    defparam full_nxt_c_I_6_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i1_2_lut_adj_38 (.I0(dc32_fifo_almost_full), .I1(DEBUG_1_c_c), 
            .I2(GND_net), .I3(GND_net), .O(FT_OE_N_420));   // src/fifo_dc_32_lut_gen.v(410[29] 422[32])
    defparam i1_2_lut_adj_38.LUT_INIT = 16'heeee;
    SB_LUT4 n12845_bdd_4_lut (.I0(n12845), .I1(\REG.mem_61_3 ), .I2(\REG.mem_60_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11128));
    defparam n12845_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3548_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_0_8 ), .O(n4931));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3548_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11455 (.I0(rd_addr_r_c[1]), .I1(n11507), 
            .I2(n11508), .I3(rd_addr_r_c[2]), .O(n13493));
    defparam rd_addr_r_1__bdd_4_lut_11455.LUT_INIT = 16'he4aa;
    SB_LUT4 n13493_bdd_4_lut (.I0(n13493), .I1(n11496), .I2(n11495), .I3(rd_addr_r_c[2]), 
            .O(n11562));
    defparam n13493_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i161_162 (.Q(\REG.mem_1_9 ), .C(FIFO_CLK_c), .D(n4833));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11460 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_8 ), 
            .I2(\REG.mem_3_8 ), .I3(rd_addr_r_c[1]), .O(n13487));
    defparam rd_addr_r_0__bdd_4_lut_11460.LUT_INIT = 16'he4aa;
    SB_LUT4 n13487_bdd_4_lut (.I0(n13487), .I1(\REG.mem_1_8 ), .I2(\REG.mem_0_8 ), 
            .I3(rd_addr_r_c[1]), .O(n13490));
    defparam n13487_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10940 (.I0(rd_addr_r_c[3]), .I1(n12746), 
            .I2(n11070), .I3(rd_addr_r_c[4]), .O(n12839));
    defparam rd_addr_r_3__bdd_4_lut_10940.LUT_INIT = 16'he4aa;
    SB_LUT4 i3549_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_0_7 ), .O(n4932));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3549_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11480 (.I0(rd_addr_r_c[3]), .I1(n11888), 
            .I2(n11889), .I3(rd_addr_r_c[4]), .O(n13481));
    defparam rd_addr_r_3__bdd_4_lut_11480.LUT_INIT = 16'he4aa;
    SB_LUT4 n13481_bdd_4_lut (.I0(n13481), .I1(n11877), .I2(n13394), .I3(rd_addr_r_c[4]), 
            .O(n13484));
    defparam n13481_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i179_180 (.Q(\REG.mem_1_15 ), .C(FIFO_CLK_c), .D(n4832));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12839_bdd_4_lut (.I0(n12839), .I1(n11025), .I2(n12692), .I3(rd_addr_r_c[4]), 
            .O(n12842));
    defparam n12839_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_en_i_I_0_2_lut (.I0(DEBUG_5_c), .I1(full_o), .I2(GND_net), 
            .I3(GND_net), .O(wr_sig_mv_w));   // src/fifo_dc_32_lut_gen.v(293[28:49])
    defparam wr_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10910 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_13 ), 
            .I2(\REG.mem_63_13 ), .I3(rd_addr_r_c[1]), .O(n12833));
    defparam rd_addr_r_0__bdd_4_lut_10910.LUT_INIT = 16'he4aa;
    SB_LUT4 n12833_bdd_4_lut (.I0(n12833), .I1(\REG.mem_61_13 ), .I2(\REG.mem_60_13 ), 
            .I3(rd_addr_r_c[1]), .O(n12836));
    defparam n12833_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11445 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_3 ), 
            .I2(\REG.mem_27_3 ), .I3(rd_addr_r_c[1]), .O(n13475));
    defparam rd_addr_r_0__bdd_4_lut_11445.LUT_INIT = 16'he4aa;
    SB_DFF i164_165 (.Q(\REG.mem_1_10 ), .C(FIFO_CLK_c), .D(n4831));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3550_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_0_6 ), .O(n4933));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3550_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i18_2_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n18_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i18_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3551_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_0_5 ), .O(n4934));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3551_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3552_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_0_4 ), .O(n4935));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3552_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13475_bdd_4_lut (.I0(n13475), .I1(\REG.mem_25_3 ), .I2(\REG.mem_24_3 ), 
            .I3(rd_addr_r_c[1]), .O(n11068));
    defparam n13475_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3557_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_0_3 ), .O(n4940));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3557_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10900 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_0 ), 
            .I2(\REG.mem_27_0 ), .I3(rd_addr_r_c[1]), .O(n12827));
    defparam rd_addr_r_0__bdd_4_lut_10900.LUT_INIT = 16'he4aa;
    SB_LUT4 i3558_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_0_2 ), .O(n4941));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3558_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12827_bdd_4_lut (.I0(n12827), .I1(\REG.mem_25_0 ), .I2(\REG.mem_24_0 ), 
            .I3(rd_addr_r_c[1]), .O(n12830));
    defparam n12827_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3560_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_0_1 ), .O(n4943));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3560_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11435 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_5 ), 
            .I2(\REG.mem_11_5 ), .I3(rd_addr_r_c[1]), .O(n13469));
    defparam rd_addr_r_0__bdd_4_lut_11435.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i38_2_lut_3_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n38));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i38_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10895 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_9 ), 
            .I2(\REG.mem_47_9 ), .I3(rd_addr_r_c[1]), .O(n12821));
    defparam rd_addr_r_0__bdd_4_lut_10895.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i102_2_lut_3_lut_4_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n49));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i102_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 n13469_bdd_4_lut (.I0(n13469), .I1(\REG.mem_9_5 ), .I2(\REG.mem_8_5 ), 
            .I3(rd_addr_r_c[1]), .O(n13472));
    defparam n13469_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12821_bdd_4_lut (.I0(n12821), .I1(\REG.mem_45_9 ), .I2(\REG.mem_44_9 ), 
            .I3(rd_addr_r_c[1]), .O(n12824));
    defparam n12821_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i101_2_lut_3_lut_4_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n17));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i101_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i116_2_lut_3_lut (.I0(n36), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n42));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i116_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i115_2_lut_3_lut (.I0(n36), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n10));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i115_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10990 (.I0(rd_addr_r_c[2]), .I1(n11464), 
            .I2(n11485), .I3(rd_addr_r_c[3]), .O(n12815));
    defparam rd_addr_r_2__bdd_4_lut_10990.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11450 (.I0(rd_addr_r_c[1]), .I1(n11915), 
            .I2(n11916), .I3(rd_addr_r_c[2]), .O(n13463));
    defparam rd_addr_r_1__bdd_4_lut_11450.LUT_INIT = 16'he4aa;
    SB_LUT4 i4079_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_33_4 ), .O(n5462));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4079_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13463_bdd_4_lut (.I0(n13463), .I1(n11892), .I2(n11891), .I3(rd_addr_r_c[2]), 
            .O(n11070));
    defparam n13463_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10504 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_2 ), 
            .I2(\REG.mem_15_2 ), .I3(rd_addr_r_c[1]), .O(n12347));
    defparam rd_addr_r_0__bdd_4_lut_10504.LUT_INIT = 16'he4aa;
    SB_LUT4 n12815_bdd_4_lut (.I0(n12815), .I1(n11407), .I2(n12374), .I3(rd_addr_r_c[3]), 
            .O(n11728));
    defparam n12815_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10890 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_1 ), 
            .I2(\REG.mem_63_1 ), .I3(rd_addr_r_c[1]), .O(n12809));
    defparam rd_addr_r_0__bdd_4_lut_10890.LUT_INIT = 16'he4aa;
    SB_LUT4 n12809_bdd_4_lut (.I0(n12809), .I1(\REG.mem_61_1 ), .I2(\REG.mem_60_1 ), 
            .I3(rd_addr_r_c[1]), .O(n12812));
    defparam n12809_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4078_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_33_3 ), .O(n5461));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4078_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11430 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_12 ), 
            .I2(\REG.mem_11_12 ), .I3(rd_addr_r_c[1]), .O(n13457));
    defparam rd_addr_r_0__bdd_4_lut_11430.LUT_INIT = 16'he4aa;
    SB_LUT4 n13457_bdd_4_lut (.I0(n13457), .I1(\REG.mem_9_12 ), .I2(\REG.mem_8_12 ), 
            .I3(rd_addr_r_c[1]), .O(n13460));
    defparam n13457_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i347_348 (.Q(\REG.mem_3_7 ), .C(FIFO_CLK_c), .D(n4968));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i344_345 (.Q(\REG.mem_3_6 ), .C(FIFO_CLK_c), .D(n4967));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9409_3_lut (.I0(\REG.mem_30_9 ), .I1(\REG.mem_31_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11247));
    defparam i9409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9408_3_lut (.I0(\REG.mem_28_9 ), .I1(\REG.mem_29_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11246));
    defparam i9408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i15_2_lut (.I0(n12_adj_33), .I1(wr_addr_r[2]), 
            .I2(GND_net), .I3(GND_net), .O(n15_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i15_2_lut.LUT_INIT = 16'h8888;
    SB_DFF i341_342 (.Q(\REG.mem_3_5 ), .C(FIFO_CLK_c), .D(n4966));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i338_339 (.Q(\REG.mem_3_4 ), .C(FIFO_CLK_c), .D(n4965));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i132_2_lut_3_lut (.I0(n35), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n34));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i132_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i335_336 (.Q(\REG.mem_3_3 ), .C(FIFO_CLK_c), .D(n4964));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11425 (.I0(rd_addr_r_c[1]), .I1(n12026), 
            .I2(n12027), .I3(rd_addr_r_c[2]), .O(n13451));
    defparam rd_addr_r_1__bdd_4_lut_11425.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10925 (.I0(rd_addr_r_c[1]), .I1(n11984), 
            .I2(n11985), .I3(rd_addr_r_c[2]), .O(n12797));
    defparam rd_addr_r_1__bdd_4_lut_10925.LUT_INIT = 16'he4aa;
    SB_LUT4 i4452_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_54_15 ), .O(n5835));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4452_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13451_bdd_4_lut (.I0(n13451), .I1(n11973), .I2(n11972), .I3(rd_addr_r_c[2]), 
            .O(n13454));
    defparam n13451_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4451_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_54_14 ), .O(n5834));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4451_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12797_bdd_4_lut (.I0(n12797), .I1(n11979), .I2(n11978), .I3(rd_addr_r_c[2]), 
            .O(n12800));
    defparam n12797_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4450_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_54_13 ), .O(n5833));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4450_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4449_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_54_12 ), .O(n5832));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4449_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4448_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_54_11 ), .O(n5831));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4448_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11420 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_8 ), 
            .I2(\REG.mem_31_8 ), .I3(rd_addr_r_c[1]), .O(n13445));
    defparam rd_addr_r_0__bdd_4_lut_11420.LUT_INIT = 16'he4aa;
    SB_LUT4 n13445_bdd_4_lut (.I0(n13445), .I1(\REG.mem_29_8 ), .I2(\REG.mem_28_8 ), 
            .I3(rd_addr_r_c[1]), .O(n13448));
    defparam n13445_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i332_333 (.Q(\REG.mem_3_2 ), .C(FIFO_CLK_c), .D(n4963));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4447_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_54_10 ), .O(n5830));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4447_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4446_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_54_9 ), .O(n5829));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4446_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4445_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_54_8 ), .O(n5828));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4445_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4077_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_33_2 ), .O(n5460));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4077_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i131_2_lut_3_lut (.I0(n35), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n2));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i131_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i4444_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_54_7 ), .O(n5827));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4444_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4443_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_54_6 ), .O(n5826));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4443_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4442_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_54_5 ), .O(n5825));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4442_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10885 (.I0(rd_addr_r_c[2]), .I1(n11044), 
            .I2(n11056), .I3(rd_addr_r_c[3]), .O(n12791));
    defparam rd_addr_r_2__bdd_4_lut_10885.LUT_INIT = 16'he4aa;
    SB_LUT4 n12791_bdd_4_lut (.I0(n12791), .I1(n11041), .I2(n11035), .I3(rd_addr_r_c[3]), 
            .O(n11131));
    defparam n12791_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4441_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_54_4 ), .O(n5824));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4441_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11410 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_1 ), 
            .I2(\REG.mem_43_1 ), .I3(rd_addr_r_c[1]), .O(n13439));
    defparam rd_addr_r_0__bdd_4_lut_11410.LUT_INIT = 16'he4aa;
    SB_LUT4 i4440_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_54_3 ), .O(n5823));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4440_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10905 (.I0(rd_addr_r_c[3]), .I1(n12020), 
            .I2(n12021), .I3(rd_addr_r_c[4]), .O(n12785));
    defparam rd_addr_r_3__bdd_4_lut_10905.LUT_INIT = 16'he4aa;
    SB_LUT4 n13439_bdd_4_lut (.I0(n13439), .I1(\REG.mem_41_1 ), .I2(\REG.mem_40_1 ), 
            .I3(rd_addr_r_c[1]), .O(n13442));
    defparam n13439_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i329_330 (.Q(\REG.mem_3_1 ), .C(FIFO_CLK_c), .D(n4962));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4439_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_54_2 ), .O(n5822));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4439_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12785_bdd_4_lut (.I0(n12785), .I1(n12003), .I2(n12002), .I3(rd_addr_r_c[4]), 
            .O(n12788));
    defparam n12785_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i326_327 (.Q(\REG.mem_3_0 ), .C(FIFO_CLK_c), .D(n4961));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12347_bdd_4_lut (.I0(n12347), .I1(\REG.mem_13_2 ), .I2(\REG.mem_12_2 ), 
            .I3(rd_addr_r_c[1]), .O(n12350));
    defparam n12347_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10880 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_12 ), 
            .I2(\REG.mem_47_12 ), .I3(rd_addr_r_c[1]), .O(n12779));
    defparam rd_addr_r_0__bdd_4_lut_10880.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i36_2_lut_3_lut (.I0(n11), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n36));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i36_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i4438_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_54_1 ), .O(n5821));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4438_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4437_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_54_0 ), .O(n5820));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4437_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i275_276 (.Q(\REG.mem_2_15 ), .C(FIFO_CLK_c), .D(n4960));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11415 (.I0(rd_addr_r_c[1]), .I1(n11465), 
            .I2(n11466), .I3(rd_addr_r_c[2]), .O(n13433));
    defparam rd_addr_r_1__bdd_4_lut_11415.LUT_INIT = 16'he4aa;
    SB_DFF i272_273 (.Q(\REG.mem_2_14 ), .C(FIFO_CLK_c), .D(n4959));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4076_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_33_1 ), .O(n5459));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4076_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i35_2_lut_3_lut (.I0(n11), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n35));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i35_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i4107_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_34_15 ), .O(n5490));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4107_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i269_270 (.Q(\REG.mem_2_13 ), .C(FIFO_CLK_c), .D(n4958));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4075_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_33_0 ), .O(n5458));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4075_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12779_bdd_4_lut (.I0(n12779), .I1(\REG.mem_45_12 ), .I2(\REG.mem_44_12 ), 
            .I3(rd_addr_r_c[1]), .O(n12782));
    defparam n12779_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i266_267 (.Q(\REG.mem_2_12 ), .C(FIFO_CLK_c), .D(n4957));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13433_bdd_4_lut (.I0(n13433), .I1(n11445), .I2(n11444), .I3(rd_addr_r_c[2]), 
            .O(n11583));
    defparam n13433_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i82_2_lut_3_lut_4_lut (.I0(n17_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n59));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i82_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_DFF i263_264 (.Q(\REG.mem_2_11 ), .C(FIFO_CLK_c), .D(n4956));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wr_addr_r_6__I_0_141_7_lut (.I0(GND_net), .I1(wr_addr_r[5]), 
            .I2(GND_net), .I3(n10137), .O(wr_addr_p1_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF i260_261 (.Q(\REG.mem_2_10 ), .C(FIFO_CLK_c), .D(n4955));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i81_2_lut_3_lut_4_lut (.I0(n17_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n27));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i81_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i4106_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_34_14 ), .O(n5489));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4106_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4436_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_53_15 ), .O(n5819));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4436_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4105_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_34_13 ), .O(n5488));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4105_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4435_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_53_14 ), .O(n5818));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4435_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4434_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_53_13 ), .O(n5817));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4434_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4433_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_53_12 ), .O(n5816));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4433_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4104_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_34_12 ), .O(n5487));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4104_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4432_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_53_11 ), .O(n5815));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4432_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4431_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_53_10 ), .O(n5814));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4431_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4103_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_34_11 ), .O(n5486));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4103_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11400 (.I0(rd_addr_r_c[1]), .I1(n11537), 
            .I2(n11538), .I3(rd_addr_r_c[2]), .O(n13427));
    defparam rd_addr_r_1__bdd_4_lut_11400.LUT_INIT = 16'he4aa;
    SB_LUT4 i4430_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_53_9 ), .O(n5813));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4430_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4429_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_53_8 ), .O(n5812));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4429_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i257_258 (.Q(\REG.mem_2_9 ), .C(FIFO_CLK_c), .D(n4954));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4102_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_34_10 ), .O(n5485));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4102_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9684_3_lut (.I0(\REG.mem_32_1 ), .I1(\REG.mem_33_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11522));
    defparam i9684_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i254_255 (.Q(\REG.mem_2_8 ), .C(FIFO_CLK_c), .D(n4953));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i17_2_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n17_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i17_2_lut.LUT_INIT = 16'h8888;
    SB_DFF i251_252 (.Q(\REG.mem_2_7 ), .C(FIFO_CLK_c), .D(n4952));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13427_bdd_4_lut (.I0(n13427), .I1(n11535), .I2(n11534), .I3(rd_addr_r_c[2]), 
            .O(n11586));
    defparam n13427_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i248_249 (.Q(\REG.mem_2_6 ), .C(FIFO_CLK_c), .D(n4951));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4428_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_53_7 ), .O(n5811));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4428_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4101_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_34_9 ), .O(n5484));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4101_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4100_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_34_8 ), .O(n5483));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4100_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11395 (.I0(rd_addr_r_c[1]), .I1(n11546), 
            .I2(n11547), .I3(rd_addr_r_c[2]), .O(n13421));
    defparam rd_addr_r_1__bdd_4_lut_11395.LUT_INIT = 16'he4aa;
    SB_LUT4 i9685_3_lut (.I0(\REG.mem_34_1 ), .I1(\REG.mem_35_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11523));
    defparam i9685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4427_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_53_6 ), .O(n5810));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4427_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4099_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_34_7 ), .O(n5482));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4099_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9574_3_lut (.I0(\REG.mem_34_7 ), .I1(\REG.mem_35_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11412));
    defparam i9574_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9573_3_lut (.I0(\REG.mem_32_7 ), .I1(\REG.mem_33_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11411));
    defparam i9573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9447_3_lut (.I0(\REG.mem_4_0 ), .I1(\REG.mem_5_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11285));
    defparam i9447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9448_3_lut (.I0(\REG.mem_6_0 ), .I1(\REG.mem_7_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11286));
    defparam i9448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4426_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_53_5 ), .O(n5809));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4426_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9445_3_lut (.I0(\REG.mem_2_0 ), .I1(\REG.mem_3_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11283));
    defparam i9445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9444_3_lut (.I0(\REG.mem_0_0 ), .I1(\REG.mem_1_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11282));
    defparam i9444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9651_3_lut (.I0(\REG.mem_36_10 ), .I1(\REG.mem_37_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11489));
    defparam i9651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9652_3_lut (.I0(\REG.mem_38_10 ), .I1(\REG.mem_39_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11490));
    defparam i9652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4425_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_53_4 ), .O(n5808));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4425_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9640_3_lut (.I0(\REG.mem_34_10 ), .I1(\REG.mem_35_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11478));
    defparam i9640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9639_3_lut (.I0(\REG.mem_32_10 ), .I1(\REG.mem_33_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11477));
    defparam i9639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9612_3_lut (.I0(\REG.mem_20_10 ), .I1(\REG.mem_21_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11450));
    defparam i9612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9613_3_lut (.I0(\REG.mem_22_10 ), .I1(\REG.mem_23_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11451));
    defparam i9613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4424_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_53_3 ), .O(n5807));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4424_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9610_3_lut (.I0(\REG.mem_18_10 ), .I1(\REG.mem_19_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11448));
    defparam i9610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9609_3_lut (.I0(\REG.mem_16_10 ), .I1(\REG.mem_17_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11447));
    defparam i9609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9405_3_lut (.I0(\REG.mem_4_7 ), .I1(\REG.mem_5_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11243));
    defparam i9405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9406_3_lut (.I0(\REG.mem_6_7 ), .I1(\REG.mem_7_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11244));
    defparam i9406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10083_3_lut (.I0(n12710), .I1(n12632), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11921));
    defparam i10083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10084_3_lut (.I0(n12512), .I1(n12410), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11922));
    defparam i10084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10063_3_lut (.I0(n12920), .I1(n12782), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11901));
    defparam i10063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10062_3_lut (.I0(n13004), .I1(n12974), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11900));
    defparam i10062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4423_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_53_2 ), .O(n5806));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4423_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9364_3_lut (.I0(\REG.mem_2_7 ), .I1(\REG.mem_3_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11202));
    defparam i9364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9363_3_lut (.I0(\REG.mem_0_7 ), .I1(\REG.mem_1_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11201));
    defparam i9363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4422_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_53_1 ), .O(n5805));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4422_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9585_3_lut (.I0(\REG.mem_4_10 ), .I1(\REG.mem_5_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11423));
    defparam i9585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9586_3_lut (.I0(\REG.mem_6_10 ), .I1(\REG.mem_7_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11424));
    defparam i9586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9577_3_lut (.I0(\REG.mem_2_10 ), .I1(\REG.mem_3_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11415));
    defparam i9577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9576_3_lut (.I0(\REG.mem_0_10 ), .I1(\REG.mem_1_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11414));
    defparam i9576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4421_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_53_0 ), .O(n5804));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4421_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9634_3_lut (.I0(n13388), .I1(n13202), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11472));
    defparam i9634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9622_3_lut (.I0(n13472), .I1(n12776), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11460));
    defparam i9622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9564_3_lut (.I0(\REG.mem_52_5 ), .I1(\REG.mem_53_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11402));
    defparam i9564_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9565_3_lut (.I0(\REG.mem_54_5 ), .I1(\REG.mem_55_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11403));
    defparam i9565_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9547_3_lut (.I0(\REG.mem_50_5 ), .I1(\REG.mem_51_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11385));
    defparam i9547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9546_3_lut (.I0(\REG.mem_48_5 ), .I1(\REG.mem_49_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11384));
    defparam i9546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i80_2_lut_3_lut_4_lut (.I0(n15_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n60));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i80_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i79_2_lut_3_lut_4_lut (.I0(n15_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n28));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i79_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i3_2_lut (.I0(\rd_addr_nxt_c_6__N_498[2] ), 
            .I1(\rd_addr_nxt_c_6__N_498[3] ), .I2(GND_net), .I3(GND_net), 
            .O(rd_grey_w[2]));   // src/fifo_dc_32_lut_gen.v(504[28:66])
    defparam rd_addr_nxt_c_6__I_0_152_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4420_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_52_15 ), .O(n5803));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4420_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10067_3_lut (.I0(n13424), .I1(n11904), .I2(rd_addr_r_c[3]), 
            .I3(GND_net), .O(n11905));
    defparam i10067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10066_3_lut (.I0(n13442), .I1(n13358), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11904));
    defparam i10066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4419_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_52_14 ), .O(n5802));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4419_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9366_3_lut (.I0(\REG.mem_20_5 ), .I1(\REG.mem_21_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11204));
    defparam i9366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9367_3_lut (.I0(\REG.mem_22_5 ), .I1(\REG.mem_23_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11205));
    defparam i9367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9325_3_lut (.I0(\REG.mem_18_5 ), .I1(\REG.mem_19_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11163));
    defparam i9325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9324_3_lut (.I0(\REG.mem_16_5 ), .I1(\REG.mem_17_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11162));
    defparam i9324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4418_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_52_13 ), .O(n5801));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4418_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4417_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_52_12 ), .O(n5800));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4417_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4416_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_52_11 ), .O(n5799));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4416_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9234_3_lut (.I0(\REG.mem_4_5 ), .I1(\REG.mem_5_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11072));
    defparam i9234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9235_3_lut (.I0(\REG.mem_6_5 ), .I1(\REG.mem_7_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11073));
    defparam i9235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4415_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_52_10 ), .O(n5798));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4415_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i47_2_lut_3_lut_4_lut (.I0(n12_adj_33), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n47_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i47_2_lut_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 EnabledDecoder_2_i49_2_lut_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n49_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i49_2_lut_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i4414_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_52_9 ), .O(n5797));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4414_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10098_3_lut (.I0(\REG.mem_60_8 ), .I1(\REG.mem_61_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11936));
    defparam i10098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10099_3_lut (.I0(\REG.mem_62_8 ), .I1(\REG.mem_63_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11937));
    defparam i10099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9199_3_lut (.I0(\REG.mem_2_5 ), .I1(\REG.mem_3_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11037));
    defparam i9199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9198_3_lut (.I0(\REG.mem_0_5 ), .I1(\REG.mem_1_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11036));
    defparam i9198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10036_3_lut (.I0(\REG.mem_58_8 ), .I1(\REG.mem_59_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11874));
    defparam i10036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10035_3_lut (.I0(\REG.mem_56_8 ), .I1(\REG.mem_57_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11873));
    defparam i10035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_5__I_0_i6_2_lut_3_lut (.I0(wr_addr_r[5]), .I1(rp_sync2_r[5]), 
            .I2(rp_sync2_r[6]), .I3(GND_net), .O(n6_adj_37));   // src/fifo_dc_32_lut_gen.v(295[31:67])
    defparam wr_addr_r_5__I_0_i6_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4413_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_52_8 ), .O(n5796));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4413_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut (.I0(rp_sync2_r[2]), .I1(rp_sync2_r[3]), .I2(rp_sync_w[4]), 
            .I3(GND_net), .O(rp_sync_w[2]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_39 (.I0(rp_sync2_r[0]), .I1(rp_sync2_r[1]), 
            .I2(rp_sync_w[2]), .I3(GND_net), .O(rp_sync_w[0]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_3_lut_adj_39.LUT_INIT = 16'h9696;
    SB_LUT4 i4098_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_34_6 ), .O(n5481));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4098_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_fifo_en_w_I_0_158_2_lut_3_lut (.I0(DEBUG_3_c), .I1(get_next_word), 
            .I2(\genblk16.rd_prev_r ), .I3(GND_net), .O(t_rd_fifo_en_w));   // src/fifo_dc_32_lut_gen.v(747[41:67])
    defparam rd_fifo_en_w_I_0_158_2_lut_3_lut.LUT_INIT = 16'hf4f4;
    SB_LUT4 i10089_3_lut (.I0(\REG.mem_60_15 ), .I1(\REG.mem_61_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11927));
    defparam i10089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10090_3_lut (.I0(\REG.mem_62_15 ), .I1(\REG.mem_63_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11928));
    defparam i10090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10081_3_lut (.I0(\REG.mem_58_15 ), .I1(\REG.mem_59_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11919));
    defparam i10081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10080_3_lut (.I0(\REG.mem_56_15 ), .I1(\REG.mem_57_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11918));
    defparam i10080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4097_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_34_5 ), .O(n5480));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4097_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4096_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_34_4 ), .O(n5479));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4096_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4412_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_52_7 ), .O(n5795));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4412_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4411_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_52_6 ), .O(n5794));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4411_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4410_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_52_5 ), .O(n5793));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4410_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4409_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_52_4 ), .O(n5792));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4409_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i57_2_lut_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n57_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i57_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i9441_3_lut (.I0(\REG.mem_36_9 ), .I1(\REG.mem_37_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11279));
    defparam i9441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9442_3_lut (.I0(\REG.mem_38_9 ), .I1(\REG.mem_39_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11280));
    defparam i9442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9415_3_lut (.I0(\REG.mem_34_9 ), .I1(\REG.mem_35_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11253));
    defparam i9415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9414_3_lut (.I0(\REG.mem_32_9 ), .I1(\REG.mem_33_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11252));
    defparam i9414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9372_3_lut (.I0(\REG.mem_20_9 ), .I1(\REG.mem_21_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11210));
    defparam i9372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9373_3_lut (.I0(\REG.mem_22_9 ), .I1(\REG.mem_23_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11211));
    defparam i9373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9349_3_lut (.I0(\REG.mem_18_9 ), .I1(\REG.mem_19_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11187));
    defparam i9349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9348_3_lut (.I0(\REG.mem_16_9 ), .I1(\REG.mem_17_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11186));
    defparam i9348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i59_2_lut_3_lut_4_lut (.I0(n11), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n59_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i59_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i9_2_lut_3_lut_4_lut (.I0(DEBUG_5_c), .I1(full_o), 
            .I2(wr_addr_r[0]), .I3(wr_addr_r[1]), .O(n9));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i9_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i4408_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_52_3 ), .O(n5791));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4408_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i42_2_lut_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n42_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i42_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i4095_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_34_3 ), .O(n5478));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4095_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4407_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_52_2 ), .O(n5790));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4407_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9051_4_lut_4_lut (.I0(rd_addr_r_c[1]), .I1(rd_addr_r_c[2]), 
            .I2(wp_sync2_r[1]), .I3(wp_sync_w[2]), .O(n10887));
    defparam i9051_4_lut_4_lut.LUT_INIT = 16'hb7de;
    SB_LUT4 i1_2_lut_3_lut_adj_40 (.I0(wp_sync2_r[4]), .I1(wp_sync2_r[6]), 
            .I2(wp_sync2_r[5]), .I3(GND_net), .O(wp_sync_w[4]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_adj_40.LUT_INIT = 16'h9696;
    SB_LUT4 i9594_3_lut (.I0(\REG.mem_60_5 ), .I1(\REG.mem_61_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11432));
    defparam i9594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9595_3_lut (.I0(\REG.mem_62_5 ), .I1(\REG.mem_63_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11433));
    defparam i9595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_41 (.I0(wp_sync2_r[0]), .I1(wp_sync2_r[1]), 
            .I2(wp_sync_w[2]), .I3(GND_net), .O(wp_sync_w[0]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_adj_41.LUT_INIT = 16'h9696;
    SB_LUT4 EnabledDecoder_2_i63_2_lut_3_lut_4_lut (.I0(n12_adj_33), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n63));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i63_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_3_lut_adj_42 (.I0(wp_sync2_r[2]), .I1(wp_sync2_r[3]), 
            .I2(wp_sync_w[4]), .I3(GND_net), .O(wp_sync_w[2]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_adj_42.LUT_INIT = 16'h9696;
    SB_LUT4 i9583_3_lut (.I0(\REG.mem_58_5 ), .I1(\REG.mem_59_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11421));
    defparam i9583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9582_3_lut (.I0(\REG.mem_56_5 ), .I1(\REG.mem_57_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11420));
    defparam i9582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4406_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_52_1 ), .O(n5789));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4406_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i65_2_lut_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n65));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i65_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i9655_3_lut (.I0(n12464), .I1(n12344), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11493));
    defparam i9655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9654_3_lut (.I0(n12890), .I1(n12584), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11492));
    defparam i9654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4405_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_52_0 ), .O(n5788));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4405_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9737_3_lut (.I0(n13058), .I1(n11574), .I2(rd_addr_r_c[3]), 
            .I3(GND_net), .O(n11575));
    defparam i9737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9736_3_lut (.I0(n12998), .I1(n12926), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11574));
    defparam i9736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10076_3_lut (.I0(n13454), .I1(n11913), .I2(rd_addr_r_c[3]), 
            .I3(GND_net), .O(n11914));
    defparam i10076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10075_3_lut (.I0(n13784), .I1(n13256), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11913));
    defparam i10075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9411_3_lut (.I0(n12302), .I1(n13664), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11249));
    defparam i9411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9396_3_lut (.I0(\REG.mem_52_4 ), .I1(\REG.mem_53_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11234));
    defparam i9396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9397_3_lut (.I0(\REG.mem_54_4 ), .I1(\REG.mem_55_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11235));
    defparam i9397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9388_3_lut (.I0(\REG.mem_50_4 ), .I1(\REG.mem_51_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11226));
    defparam i9388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9387_3_lut (.I0(\REG.mem_48_4 ), .I1(\REG.mem_49_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11225));
    defparam i9387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9375_3_lut (.I0(\REG.mem_36_4 ), .I1(\REG.mem_37_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11213));
    defparam i9375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9376_3_lut (.I0(\REG.mem_38_4 ), .I1(\REG.mem_39_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11214));
    defparam i9376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9370_3_lut (.I0(\REG.mem_34_4 ), .I1(\REG.mem_35_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11208));
    defparam i9370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9369_3_lut (.I0(\REG.mem_32_4 ), .I1(\REG.mem_33_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11207));
    defparam i9369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9351_3_lut (.I0(\REG.mem_20_4 ), .I1(\REG.mem_21_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11189));
    defparam i9351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9352_3_lut (.I0(\REG.mem_22_4 ), .I1(\REG.mem_23_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11190));
    defparam i9352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9340_3_lut (.I0(\REG.mem_18_4 ), .I1(\REG.mem_19_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11178));
    defparam i9340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9339_3_lut (.I0(\REG.mem_16_4 ), .I1(\REG.mem_17_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11177));
    defparam i9339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9190_3_lut (.I0(n12392), .I1(n12356), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11028));
    defparam i9190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9189_3_lut (.I0(n12626), .I1(n12530), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11027));
    defparam i9189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9597_3_lut (.I0(\REG.mem_12_10 ), .I1(\REG.mem_13_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11435));
    defparam i9597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9598_3_lut (.I0(\REG.mem_14_10 ), .I1(\REG.mem_15_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11436));
    defparam i9598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9589_3_lut (.I0(\REG.mem_10_10 ), .I1(\REG.mem_11_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11427));
    defparam i9589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9588_3_lut (.I0(\REG.mem_8_10 ), .I1(\REG.mem_9_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11426));
    defparam i9588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i45_2_lut_3_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n45));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i45_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i78_2_lut_3_lut_4_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n61));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i78_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i77_2_lut_3_lut_4_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n29));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i77_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i4404_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_51_15 ), .O(n5787));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4404_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4403_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_51_14 ), .O(n5786));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4403_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4402_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_51_13 ), .O(n5785));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4402_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4401_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_51_12 ), .O(n5784));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4401_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4400_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_51_11 ), .O(n5783));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4400_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9630_3_lut (.I0(\REG.mem_28_10 ), .I1(\REG.mem_29_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11468));
    defparam i9630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9631_3_lut (.I0(\REG.mem_30_10 ), .I1(\REG.mem_31_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11469));
    defparam i9631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4399_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_51_10 ), .O(n5782));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4399_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4398_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_51_9 ), .O(n5781));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4398_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4397_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_51_8 ), .O(n5780));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4397_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4396_3_lut_4_lut (.I0(n43), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_51_7 ), .O(n5779));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4396_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9619_3_lut (.I0(\REG.mem_26_10 ), .I1(\REG.mem_27_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11457));
    defparam i9619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9618_3_lut (.I0(\REG.mem_24_10 ), .I1(\REG.mem_25_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11456));
    defparam i9618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9669_3_lut (.I0(\REG.mem_44_10 ), .I1(\REG.mem_45_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11507));
    defparam i9669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9670_3_lut (.I0(\REG.mem_46_10 ), .I1(\REG.mem_47_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11508));
    defparam i9670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9658_3_lut (.I0(\REG.mem_42_10 ), .I1(\REG.mem_43_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11496));
    defparam i9658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9657_3_lut (.I0(\REG.mem_40_10 ), .I1(\REG.mem_41_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11495));
    defparam i9657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10050_3_lut (.I0(n13322), .I1(n13262), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11888));
    defparam i10050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10051_3_lut (.I0(n13196), .I1(n13130), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11889));
    defparam i10051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10039_3_lut (.I0(n13460), .I1(n13382), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11877));
    defparam i10039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10077_3_lut (.I0(\REG.mem_28_14 ), .I1(\REG.mem_29_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11915));
    defparam i10077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10078_3_lut (.I0(\REG.mem_30_14 ), .I1(\REG.mem_31_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11916));
    defparam i10078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10054_3_lut (.I0(\REG.mem_26_14 ), .I1(\REG.mem_27_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11892));
    defparam i10054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10053_3_lut (.I0(\REG.mem_24_14 ), .I1(\REG.mem_25_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11891));
    defparam i10053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10188_3_lut (.I0(\REG.mem_20_13 ), .I1(\REG.mem_21_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12026));
    defparam i10188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10189_3_lut (.I0(\REG.mem_22_13 ), .I1(\REG.mem_23_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12027));
    defparam i10189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10146_3_lut (.I0(\REG.mem_36_14 ), .I1(\REG.mem_37_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11984));
    defparam i10146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10147_3_lut (.I0(\REG.mem_38_14 ), .I1(\REG.mem_39_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11985));
    defparam i10147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10135_3_lut (.I0(\REG.mem_18_13 ), .I1(\REG.mem_19_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11973));
    defparam i10135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10134_3_lut (.I0(\REG.mem_16_13 ), .I1(\REG.mem_17_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11972));
    defparam i10134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10141_3_lut (.I0(\REG.mem_34_14 ), .I1(\REG.mem_35_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11979));
    defparam i10141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10140_3_lut (.I0(\REG.mem_32_14 ), .I1(\REG.mem_33_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11978));
    defparam i10140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10183_3_lut (.I0(n13622), .I1(n13448), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n12021));
    defparam i10183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10165_3_lut (.I0(n13604), .I1(n12704), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n12003));
    defparam i10165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10164_3_lut (.I0(n13490), .I1(n13658), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n12002));
    defparam i10164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9627_3_lut (.I0(\REG.mem_44_7 ), .I1(\REG.mem_45_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11465));
    defparam i9627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9628_3_lut (.I0(\REG.mem_46_7 ), .I1(\REG.mem_47_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11466));
    defparam i9628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9607_3_lut (.I0(\REG.mem_42_7 ), .I1(\REG.mem_43_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11445));
    defparam i9607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9606_3_lut (.I0(\REG.mem_40_7 ), .I1(\REG.mem_41_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11444));
    defparam i9606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i11_2_lut_3_lut_4_lut (.I0(DEBUG_5_c), .I1(full_o), 
            .I2(wr_addr_r[0]), .I3(wr_addr_r[1]), .O(n11));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i9699_3_lut (.I0(\REG.mem_60_10 ), .I1(\REG.mem_61_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11537));
    defparam i9699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9700_3_lut (.I0(\REG.mem_62_10 ), .I1(\REG.mem_63_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11538));
    defparam i9700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i12_2_lut_3_lut_4_lut (.I0(DEBUG_5_c), .I1(full_o), 
            .I2(wr_addr_r[0]), .I3(wr_addr_r[1]), .O(n12_adj_33));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i12_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i9697_3_lut (.I0(\REG.mem_58_10 ), .I1(\REG.mem_59_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11535));
    defparam i9697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9696_3_lut (.I0(\REG.mem_56_10 ), .I1(\REG.mem_57_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11534));
    defparam i9696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i43_2_lut_3_lut_4_lut (.I0(n11), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n43));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i43_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i9708_3_lut (.I0(\REG.mem_36_1 ), .I1(\REG.mem_37_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11546));
    defparam i9708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9709_3_lut (.I0(\REG.mem_38_1 ), .I1(\REG.mem_39_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11547));
    defparam i9709_3_lut.LUT_INIT = 16'hcaca;
=======
    wire n25_c;
    wire [5:0]wr_addr_r;   // src/fifo_dc_32_lut_gen.v(196[29:38])
    
    wire \REG.mem_18_22 , n6196, \REG.mem_18_21 , n6195, \REG.mem_0_9 ;
    wire [5:0]rd_addr_r;   // src/fifo_dc_32_lut_gen.v(217[29:38])
    
    wire n13237, \REG.mem_2_9 , \REG.mem_3_9 , n13238, \REG.mem_18_20 , 
        n6194, n14647, n13064, n13063, n14650, \REG.mem_18_19 , 
        n6193, \REG.mem_18_18 , n6192, \REG.mem_18_17 , n6191, n13244, 
        n13243, \REG.mem_18_16 , n6190, n13270, \REG.mem_18_25 , \REG.mem_19_25 , 
        n15793, n14515, \REG.mem_0_31 , n14518, n15073, n14016, 
        n13271;
    wire [5:0]n1;
    
    wire \REG.mem_16_25 , n13794, \REG.mem_18_15 , n6189, n15787, 
        \REG.mem_0_7 , n13588, \REG.mem_2_7 , \REG.mem_3_7 , n13589, 
        \REG.mem_18_14 , n6188, n8_c, n13241, n13240, \REG.mem_30_9 , 
        \REG.mem_31_9 , n13277, n14641, \REG.mem_18_13 , n6187, n13812, 
        \REG.mem_28_9 , \REG.mem_29_9 , n13276, n14194, n14195, n15067, 
        \REG.mem_18_12 , n6186, \REG.mem_16_7 , n13273, \REG.mem_18_7 , 
        \REG.mem_19_7 , n13274, n13898, n13897, n14189, n14188, 
        n13157, n14644, \REG.mem_18_11 , n6185, n5704, \REG.mem_3_10 , 
        n13929, n13938, n15061, \REG.mem_18_10 , n6184, n13911, 
        n13890, n15064, \afull_flag_impl.af_flag_nxt_w , n12_c, \REG.mem_18_9 , 
        n6183, n13_c, \REG.mem_18_8 , n6182, n5703, n30, \REG.mem_29_31 , 
        n6557, n6181, \REG.mem_29_30 , n6556, n15775, \REG.mem_18_6 , 
        n6180, n13366, n13367, n15055, n15778, \REG.mem_29_29 , 
        n6555, n5702, \REG.mem_3_8 , \REG.mem_18_5 , n6179, \REG.mem_18_4 , 
        n6178, n13361, n13360, n13483, \REG.mem_14_11 , \REG.mem_15_11 , 
        n15769;
    wire [31:0]rd_data_o_31__N_598;
    
    wire rd_fifo_en_w, \REG.mem_29_28 , n6554, n15049, \REG.mem_29_27 , 
        n6553, \REG.mem_13_11 , \REG.mem_12_11 , n15772, n15763, \REG.mem_18_3 , 
        n6177, n13827, n15052, \REG.mem_0_10 , n13288, \REG.mem_2_10 , 
        n13289, \REG.mem_18_2 , n6176, \REG.mem_18_1 , n6175, \REG.mem_29_26 , 
        n6552, \REG.mem_18_0 , n6174, n13295, n13294, \REG.mem_2_26 , 
        \REG.mem_3_26 , n15043, \REG.mem_0_26 , n15046, \REG.mem_14_16 , 
        \REG.mem_15_16 , n15757, \REG.mem_29_25 , n6551, n13944, n13956, 
        n15037, n13935, n13923, n15040, \REG.mem_13_16 , \REG.mem_12_16 , 
        n13830, \REG.mem_14_5 , \REG.mem_15_5 , n15031, \REG.mem_13_5 , 
        \REG.mem_12_5 , n14025, n13309, n13310, n15751, n13292, 
        n13291, n13837, n5701, n13986, n13995, n15025, n5700, 
        \REG.mem_3_6 , n13971, n13953, n15028, n14, \REG.mem_14_29 , 
        \REG.mem_15_29 , n15745, \REG.mem_29_24 , n6550, \REG.mem_29_23 , 
        n6549, \REG.mem_13_29 , \REG.mem_12_29 , n15748, n5699, \REG.mem_3_5 ;
    wire [5:0]rd_grey_w;   // src/fifo_dc_32_lut_gen.v(224[38:47])
    
    wire n13114, n13115, n15019, empty_nxt_c_N_636;
    wire [5:0]wr_grey_w;   // src/fifo_dc_32_lut_gen.v(203[38:47])
    
    wire n5698, \REG.mem_3_4 , \REG.mem_29_22 , n6548, \REG.mem_2_31 , 
        \REG.mem_3_31 , \REG.mem_29_21 , n6547, \REG.mem_29_20 , n6546, 
        n13085, n13084, n15022, n15, \REG.mem_29_19 , n6545, n13060, 
        n13061, n15721, n14998, n13436, n15013, n13322, n13321, 
        n13838, n13729, n13730, n15715, n13694, n15496, n13433, 
        n14992, n13357, n13358, n15709, \REG.mem_29_18 , n6544, 
        n13402, n13403, n15007, n13397, n13396, n13444, \REG.mem_29_17 , 
        n6543, \REG.mem_29_16 , n6542, \REG.mem_29_15 , n6541, \REG.mem_29_14 , 
        n6540, \REG.mem_29_13 , n6539, \REG.mem_29_12 , n6538, n13738, 
        n13739, n14995, n5697, \REG.mem_3_3 , n13349, n13348, n13379, 
        n14174, n14173, \REG.mem_29_11 , n6537, \REG.mem_29_10 , n6536, 
        n6535, n14122, n14123, n14989, \REG.mem_29_8 , n6534, \REG.mem_30_25 , 
        \REG.mem_31_25 , n15691, n5696, \REG.mem_3_2 , n14566, n13690, 
        \REG.mem_28_25 , n13851, \REG.mem_29_7 , n6533, n13769, n13768, 
        n13372, n13373, n15685, n15862, n15598, n13058, \REG.mem_16_10 , 
        n13306, \REG.mem_19_10 , n13307, n13313, n13312, n7_adj_1372, 
        n8_adj_1373, n12209;
    wire [5:0]rp_sync2_r;   // src/fifo_dc_32_lut_gen.v(202[37:47])
    wire [5:0]n1_adj_1394;
    
    wire \REG.mem_29_6 , n6532, n27_c, n14902, n15640, n13852, n13364, 
        n13363, n13391, n15202, n16180, n13853, n13445, n14977, 
        \REG.mem_29_5 , n6531, \REG.mem_29_4 , n6530, \REG.mem_29_3 , 
        n6529, \REG.mem_29_2 , n6528, \REG.mem_3_1 , n5695, \REG.mem_29_1 , 
        n6527, n13418, n14968, \REG.mem_3_0 , n5694, n5725, \REG.mem_3_30 , 
        n5724, \REG.mem_3_29 , n5723, \REG.mem_29_0 , n6526, full_nxt_c_N_633, 
        \REG.mem_3_28 , n5722, n14704, n14692, n14971, n15673, \REG.mem_3_27 , 
        n5721, n14722, n14764, n14974, n5720, n15676, \REG.mem_3_25 , 
        n5719, \REG.mem_3_24 , n5718, \REG.mem_3_23 , n5717, \REG.mem_3_22 , 
        n5716, \REG.mem_3_21 , n5715, \REG.mem_14_1 , \REG.mem_15_1 , 
        n15667, \REG.mem_18_29 , \REG.mem_19_29 , n14629, \REG.mem_16_29 , 
        n14632, n5693, \REG.mem_3_20 , n5714, n28_adj_1375, \REG.mem_3_19 , 
        n5713, \REG.mem_13_1 , \REG.mem_12_1 , n15670, n13492, n13493, 
        n14623, n13387, n13388, n14965, n13481, n13480, n14626, 
        \REG.mem_3_18 , n5712, \REG.mem_3_17 , n5711, \REG.mem_3_16 , 
        n5710, \REG.mem_3_15 , n5709, \REG.mem_3_14 , n5708, \REG.mem_3_13 , 
        n5707, \REG.mem_3_12 , n5706;
    wire [5:0]rd_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(221[30:42])
    
    wire \REG.mem_3_11 , n5705, n7001, n10_c, \REG.mem_0_28 , n13786, 
        \REG.mem_2_28 , n13787, n13796, n13795, \REG.mem_0_2 , n13339, 
        \REG.mem_2_2 , n13340, n13343, n13342, \REG.mem_0_22 , n13087, 
        \REG.mem_2_22 , n13088, n13145, n13144, n15520, n15406, 
        n13685, n14878, n16132, n13741, \REG.mem_16_22 , n13351, 
        \REG.mem_19_22 , n13352, n13355, n13354, n6999, \REG.mem_18_23 , 
        \REG.mem_19_23 , n14533, n13385, n13384, n14521, n14524, 
        n14617, n32_adj_1376, \REG.mem_14_31 , n6077, n15655, n14956, 
        n14959, n15658, n13382, n14944, n14620, \REG.mem_2_21 , 
        n15649, \REG.mem_0_21 , n15652;
    wire [5:0]wp_sync2_r;   // src/fifo_dc_32_lut_gen.v(223[37:47])
    
    wire \REG.mem_2_13 , n15643, \REG.mem_0_13 , n13869, n6931, n6929, 
        n6927, n15637, n6621, \REG.mem_31_31 , n6620, \REG.mem_31_30 , 
        n6619, \REG.mem_31_29 , n6618, \REG.mem_31_28 , n6617, \REG.mem_31_27 , 
        n6616, \REG.mem_31_26 , n6615, n6614, \REG.mem_31_24 , n6613, 
        \REG.mem_31_23 , n6612, \REG.mem_31_22 , n6611, \REG.mem_31_21 , 
        n6610, \REG.mem_31_20 , n6609, \REG.mem_31_19 , n6608, \REG.mem_31_18 , 
        n6607, \REG.mem_31_17 , n6606, \REG.mem_31_16 , n6605, \REG.mem_31_15 , 
        n6604, \REG.mem_31_14 , n6603, \REG.mem_31_13 , n6602, \REG.mem_31_12 , 
        n6601, \REG.mem_31_11 , n6600, \REG.mem_31_10 , n6599, n6598, 
        \REG.mem_31_8 , n6597, \REG.mem_31_7 , n6596, \REG.mem_31_6 , 
        n6595, \REG.mem_31_5 , n6594, \REG.mem_31_4 , n6593, \REG.mem_31_3 , 
        n6592, \REG.mem_31_2 , n6591, \REG.mem_31_1 , n6590, \REG.mem_31_0 , 
        n6589, \REG.mem_30_31 , n6588, \REG.mem_30_30 , n6587, \REG.mem_30_29 , 
        n6586, \REG.mem_30_28 , n6585, \REG.mem_30_27 , n6584, \REG.mem_30_26 , 
        n6583, n6582, \REG.mem_30_24 , n6581, \REG.mem_30_23 , n6580, 
        \REG.mem_30_22 , n6579, \REG.mem_30_21 , n6578, \REG.mem_30_20 , 
        n6577, \REG.mem_30_19 , n6576, \REG.mem_30_18 , n6575, \REG.mem_30_17 , 
        n6574, \REG.mem_30_16 , n6573, \REG.mem_30_15 , n6572, \REG.mem_30_14 , 
        n6571, \REG.mem_30_13 , n6570, \REG.mem_30_12 , n6569, \REG.mem_30_11 , 
        n6568, \REG.mem_30_10 , n6567, n6566, \REG.mem_30_8 , n6565, 
        \REG.mem_30_7 , n6564, \REG.mem_30_6 , n6563, \REG.mem_30_5 , 
        n6562, \REG.mem_30_4 , n6561, \REG.mem_30_3 , n6560, \REG.mem_30_2 , 
        n6559, \REG.mem_30_1 , n6558, \REG.mem_30_0 , n6525, \REG.mem_28_31 , 
        n6524, \REG.mem_28_30 , n6523, \REG.mem_28_29 , n6522, \REG.mem_28_28 , 
        n6521, \REG.mem_28_27 , n6520, \REG.mem_28_26 , n6519, n6518, 
        \REG.mem_28_24 , n6517, \REG.mem_28_23 , n6516, \REG.mem_28_22 , 
        n6515, \REG.mem_28_21 , n6514, \REG.mem_28_20 , n6513, \REG.mem_28_19 , 
        n6512, \REG.mem_28_18 , n6511, \REG.mem_28_17 , n6510, \REG.mem_28_16 , 
        n6509, \REG.mem_28_15 , n6508, \REG.mem_28_14 , n6507, \REG.mem_28_13 , 
        n6506, \REG.mem_28_12 , n6505, \REG.mem_28_11 , n6504, \REG.mem_28_10 , 
        n6503, n6502, \REG.mem_28_8 , n6501, \REG.mem_28_7 , n6500, 
        \REG.mem_28_6 , n6499, \REG.mem_28_5 , n6498, \REG.mem_28_4 , 
        n6497, \REG.mem_28_3 , n6496, \REG.mem_28_2 , n6495, \REG.mem_28_1 , 
        n6494, \REG.mem_28_0 , n6237, \REG.mem_19_31 , n6236, \REG.mem_19_30 , 
        n6235, n6234, \REG.mem_19_28 , n6233, \REG.mem_19_27 , n6232, 
        \REG.mem_19_26 , n6231, n6230, \REG.mem_19_24 , n6229, n6228, 
        n6227, \REG.mem_19_21 , n6226, \REG.mem_19_20 , n6225, \REG.mem_19_19 , 
        n6224, \REG.mem_19_18 , n6223, \REG.mem_19_17 , n6222, \REG.mem_19_16 , 
        n6221, \REG.mem_19_15 , n6220, \REG.mem_19_14 , n6219, \REG.mem_19_13 , 
        n6218, \REG.mem_19_12 , n6217, \REG.mem_19_11 , n6216, n6215, 
        \REG.mem_19_9 , n6214, \REG.mem_19_8 , n6213, n6212, \REG.mem_19_6 , 
        n6211, \REG.mem_19_5 , n6210, \REG.mem_19_4 , n6209, \REG.mem_19_3 , 
        n6208, \REG.mem_19_2 , n6207, \REG.mem_19_1 , n6206, \REG.mem_19_0 , 
        n6205, \REG.mem_18_31 , n6204, \REG.mem_18_30 , n6203, n6202, 
        \REG.mem_18_28 , n6201, \REG.mem_18_27 , n6200, \REG.mem_18_26 , 
        n6199, n6198, \REG.mem_18_24 , n6197, n6141, \REG.mem_16_31 , 
        n6140, \REG.mem_16_30 , n6139, n6138, \REG.mem_16_28 , n6137, 
        \REG.mem_16_27 , n6136, \REG.mem_16_26 , n6135, n6134, \REG.mem_16_24 , 
        n6133, \REG.mem_16_23 , n6132, n6131, \REG.mem_16_21 , n6130, 
        \REG.mem_16_20 , n6129, \REG.mem_16_19 , n6128, \REG.mem_16_18 , 
        n6127, \REG.mem_16_17 , n6126, \REG.mem_16_16 , n6125, \REG.mem_16_15 , 
        n6124, \REG.mem_16_14 , n6123, \REG.mem_16_13 , n6122, \REG.mem_16_12 , 
        n6121, \REG.mem_16_11 , n6120, n6119, \REG.mem_16_9 , n6118, 
        \REG.mem_16_8 , n6117, n6116, \REG.mem_16_6 , n6115, \REG.mem_16_5 , 
        n6114, \REG.mem_16_4 , n6113, \REG.mem_16_3 , n6112, \REG.mem_16_2 , 
        n6111, \REG.mem_16_1 , n6110, \REG.mem_16_0 , n6109, \REG.mem_15_31 , 
        n6108, \REG.mem_15_30 , n6107, n6106, \REG.mem_15_28 , n6105, 
        \REG.mem_15_27 , n6104, \REG.mem_15_26 , n6103, \REG.mem_15_25 , 
        n6102, \REG.mem_15_24 , n6101, \REG.mem_15_23 , n6100, \REG.mem_15_22 , 
        n6099, \REG.mem_15_21 , n6098, \REG.mem_15_20 , n6097, \REG.mem_15_19 , 
        n6096, \REG.mem_15_18 , n6095, \REG.mem_15_17 , n6094, n6093, 
        \REG.mem_15_15 , n6092, \REG.mem_15_14 , n6091, \REG.mem_15_13 , 
        n6090, \REG.mem_15_12 , n6089, n6088, \REG.mem_15_10 , \REG.mem_14_30 , 
        n6076, n6087, \REG.mem_15_9 , n6086, \REG.mem_15_8 , n6085, 
        \REG.mem_15_7 , n6084, \REG.mem_15_6 , n6083, n6082, \REG.mem_15_4 , 
        n6081, \REG.mem_15_3 , n6080, \REG.mem_15_2 , n6079, n6078, 
        \REG.mem_15_0 , n14953, n6075, n6074, \REG.mem_14_28 , n6073, 
        \REG.mem_14_27 , n6072, \REG.mem_14_26 , n6071, \REG.mem_14_25 , 
        n6070, \REG.mem_14_24 , n5692, \REG.mem_2_30 , n13484, n14947, 
        n14938, n5691, \REG.mem_2_29 , n13742, n15631, n5690, n15472, 
        n14941, n14935, n6069, \REG.mem_14_23 , n14548, n15808, 
        n6068, \REG.mem_14_22 , n6067, \REG.mem_14_21 , n6066, \REG.mem_14_20 , 
        n6065, \REG.mem_14_19 , n6064, \REG.mem_14_18 , n6063, \REG.mem_14_17 , 
        n6062, n6061, \REG.mem_14_15 , n5689, \REG.mem_2_27 , \REG.mem_0_1 , 
        \REG.mem_2_1 , n5688, n14800, n14929, n5687, \REG.mem_2_25 , 
        n6060, \REG.mem_14_14 , n15625, n15628, n13139, n14746, 
        n14611, n6059, \REG.mem_14_13 , n6058, \REG.mem_14_12 , n6057, 
        n6056, \REG.mem_14_10 , n6055, \REG.mem_14_9 , n6054, \REG.mem_14_8 , 
        n6053, \REG.mem_14_7 , n14614, n5686, \REG.mem_2_24 , n5685, 
        \REG.mem_2_23 , n6052, \REG.mem_14_6 , n6051, n6050, \REG.mem_14_4 , 
        n6049, \REG.mem_14_3 , n6048, \REG.mem_14_2 , n6047, n6046, 
        \REG.mem_14_0 , n6045, \REG.mem_13_31 , n6044, \REG.mem_13_30 , 
        n15613, n15616, n14923, n13764, n13668, n15607, n6043, 
        n13761, n13683, n15610, n6042, \REG.mem_13_28 , n14926, 
        n6041, \REG.mem_13_27 , n6040, \REG.mem_13_26 , n6039, \REG.mem_13_25 , 
        n6038, \REG.mem_13_24 , n6037, \REG.mem_13_23 , n6036, \REG.mem_13_22 , 
        n6035, \REG.mem_13_21 , n6034, \REG.mem_13_20 , n6033, \REG.mem_13_19 , 
        n6032, \REG.mem_13_18 , n6031, \REG.mem_13_17 , n6030, n6029, 
        \REG.mem_13_15 , n6028, \REG.mem_13_14 , n6027, \REG.mem_13_13 , 
        n6026, \REG.mem_13_12 , n13989, n13614, n14917, n6025, n6024, 
        \REG.mem_13_10 , n6023, \REG.mem_13_9 , n6022, \REG.mem_13_8 , 
        n6021, \REG.mem_13_7 , n5684, n6020, \REG.mem_13_6 , n6019, 
        n6018, \REG.mem_13_4 , n15601, \REG.mem_12_28 , n15604, n13983, 
        n13629, n14920, n6017, \REG.mem_13_3 , n14911, n6016, \REG.mem_13_2 , 
        n5683, n6015, n5682, \REG.mem_2_20 , n14914, n15595, n6014, 
        \REG.mem_13_0 , n5681, \REG.mem_2_19 , n6013, \REG.mem_12_31 ;
    wire [5:0]rp_sync_w;   // src/fifo_dc_32_lut_gen.v(205[30:39])
    
    wire n6012, \REG.mem_12_30 , n6011, n14899, n6010, \REG.mem_0_30 , 
        n5680, \REG.mem_2_18 , n14893, n15583, n14599, \REG.mem_0_19 , 
        n13161, n21, \REG.mem_0_4 , n5562, n5679, \REG.mem_2_17 , 
        n6009, \REG.mem_12_27 , n6008, \REG.mem_12_26 , n14887, n13164, 
        n15586;
    wire [5:0]wr_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(200[30:42])
    
    wire n8_adj_1377, n5678, \REG.mem_2_16 , n12994, n14602, n12970, 
        n15571, n14794, n13154, n14881, n5677, \REG.mem_2_15 , n12958, 
        n5676, \REG.mem_2_14 , n13884, n12932, n5675, n14875, n15565, 
        n5674, \REG.mem_2_12 , n5673, \REG.mem_2_11 , n14239, n13887, 
        n13050, n12106, n14869, n14503, n14506, n14539, n14527, 
        n13650, n14530, n14497, n14500, n5584, n14872, n13325, 
        n13324, n15514, n13706, n15553, n13691, n14863, n5672, 
        n15220, n12105, n6_adj_1378, n12136, n13167, \REG.mem_2_6 , 
        n15547, n5671, n5670, \REG.mem_2_8 , n6007, \REG.mem_12_25 , 
        n6006, \REG.mem_12_24 , n6005, \REG.mem_12_23 , n6004, \REG.mem_12_22 , 
        n6003, \REG.mem_12_21 , n5669, n14593, \REG.mem_0_27 , \REG.mem_0_6 , 
        n14857, n14848, n13316, n14851, n15541, n12135, n12134, 
        n12133, n12104;
    wire [5:0]wr_sig_diff0_w;   // src/fifo_dc_32_lut_gen.v(212[30:44])
    
    wire n12103, n12132, n14596, n5668, n13304, n14842, n5667, 
        \REG.mem_2_5 , n5666, \REG.mem_2_4 , n14491, n15544, n12131, 
        n12130, n12129, n12128, n12102, n8993, n14845, n15535;
    wire [5:0]wr_addr_nxt_c;   // src/fifo_dc_32_lut_gen.v(198[29:42])
    
    wire n14839, n12127, n6_adj_1379, n12070;
    wire [5:0]rd_sig_diff0_w;   // src/fifo_dc_32_lut_gen.v(233[30:44])
    
    wire n13892, \REG.mem_2_0 , n15529, n13891, n14833, \REG.mem_0_0 , 
        n13425, n13280, n14824, n15523, n14818, n13268, n14827, 
        n13247, n14812, n14821, n13662, n15526, n5650, \REG.mem_2_3 , 
        n5649, n5642, n5641, \REG.mem_0_11 , n6002, \REG.mem_12_20 , 
        n15517, \REG.mem_0_24 , n5622, n6001, \REG.mem_12_19 , n6000, 
        \REG.mem_12_18 , n5999, \REG.mem_12_17 , n5998, n5640, n13228, 
        n13229, n14815, n13226, n13225, n13633, n13634, n15511, 
        n13216, n13217, n14809, n13712, n13711, n13214, n13213, 
        n13963, n13964, n14803, n5569, n13211, n13210, n13546, 
        n13547, n14797, n13747, n13748, n15505, n14135, n14134, 
        n14162, n14161, n5639, \REG.mem_0_12 , n5638, n5637, \REG.mem_0_14 , 
        n5634, \REG.mem_0_15 , n5633, \REG.mem_0_16 , n5632, \REG.mem_0_17 , 
        n5631, n5630, \REG.mem_0_18 , n5629, n13336, n13337, n15493, 
        n13844, n13843, n15487, \REG.mem_12_13 , n13902, n13108, 
        n13109, n14791, n13097, n13096, n5628, \REG.mem_0_20 , n14785, 
        n14788, n15481, n14779, n14782, n15484, n5997, \REG.mem_12_15 , 
        n14773, n13170;
    wire [5:0]wp_sync_w;   // src/fifo_dc_32_lut_gen.v(226[30:39])
    
    wire n12069, n46, n12068, n5996, \REG.mem_12_14 , n12067, n5995, 
        n5994, \REG.mem_12_12 , n5993, n5992, \REG.mem_12_10 , n5627, 
        n12066, n49, n5626, n5991, \REG.mem_12_9 , n5990, \REG.mem_12_8 , 
        n5989, \REG.mem_12_7 , n14767, n14770, n5988, \REG.mem_12_6 , 
        n13735, n13736, n15469, n14761, n14755, \REG.mem_12_2 , 
        n14180, n14179, n14758, n5625, n5987, n15463, n5986, \REG.mem_12_4 , 
        n5985, \REG.mem_12_3 , n5984, n5983, n5982, \REG.mem_12_0 , 
        n5624, n14749, n5623, \REG.mem_0_23 , n15466, n14752, n5621, 
        \REG.mem_0_25 , n5620, n14137, n14138, n14743, n14155, n14156, 
        n15457, n14132, n14131, n14144, n14143, n14725, n14728, 
        n14536, n14719, n15445, n14713, n13767, n15439, n13914, 
        n14716, n13974, n13998, n14707, n13632, n13926, n14710, 
        n14701, n15427, n13917, n15421, n13980, n14004, n14695, 
        n16225, n16228, n13920, n15094, n16219, n13947, n14698, 
        n15274, n16222, n16060, n15244, n15415, n14689, n16213, 
        n16216, n16207, n16210, n14683, n5617, n15403, n14013, 
        n14007, n14686, n14662, n13124, n14677, n13121, n5616, 
        n5614, \REG.mem_0_29 , n16195, n16198, n13464, n13479, n14671, 
        n15397, n14581, n13452, n14674, n16189, n16192, n14665, 
        n14668, n13099, n13100, n14659, n15391, n13091, n13090, 
        n14116, n14117, n16183, n14111, n14110, n13568, n14653, 
        n5612, n16177, n14656, n13069, n13070, n13411, n13412, 
        n15385, n16171, n16174, n13406, n13405, n13609, n13610, 
        n15379, n13604, n15346, n4814, n5613, n16153, n14545, 
        n15226, n15322, n16156, n16147, n15367, n13932, n12960, 
        n8_adj_1387, n7_adj_1388, n16150, n14584, n9_c, n13552, 
        n13553, n16141, n13544, n13543, n13583, n13654, n13655, 
        n15361, n10_adj_1389, n12277, n13016, n13799, n13798, n15364, 
        n14125, n14126, n16135, n14120, n14119, n14159, n16129, 
        n15355, n15349, n16111, n13717, n13718, n15343, n13439, 
        n13438, n16114, n13195, n13196, n16105, n13193, n13192, 
        n15337, n16099, n15340, n16102, n15331, n13576, n13577, 
        n16087, n15325, n13550, n13549, n15319, n16075, n15313, 
        n14575, n13135, n13136, n15307, n13127, n13126, n13454, 
        n15301, n16057, n13641, n15304, n5601, n15295, n16051, 
        n15289, n14578, n16039, n13054, n13055, n15277, n13582, 
        n13103, n13104, n15271, n13207, n13208, n15265, n16027, 
        n13205, n13204, n16030, n15253, n13222, n13223, n16021, 
        n15247, n15241, n34, n13220, n13219, n15235, n16015, n16018, 
        n16009, n15238, n16003, n15229, n15223, n15997, n5570, 
        n16000, n15991, n14226, n15217, n15979, n14229, n15973, 
        n14232, n15967, n15205, n15199, n15961, n15955, n14235, 
        n15187, n13234, n13235, n15949, n13232, n13231, n15181, 
        n15184, n15943, n13594, n13595, n15937, n15175, n13562, 
        n13561, n13255, n13256, n15931, n15169, n13250, n13249, 
        n14215, n14216, n15163, n14213, n14212, n15166, n15151, 
        n14158, n15913, n14141, n14140, n13696, n13697, n15907, 
        n13643, n13642, n13567, n15901, n14494, n14129, n14128, 
        n15145, n13261, n13262, n15895, n13253, n13252, n15139, 
        n14563, n13201, n13202, n15889, n13199, n13198, n13111, 
        n13112, n15883, n14557, n13106, n13105, n13624, n13625, 
        n15877, n13592, n13591, n13285, n13286, n15871, n13283, 
        n13282, n15127, n13657, n13658, n15865, n5579, \REG.mem_0_8 , 
        n14560, n5568, \REG.mem_0_5 , n13616, n13615, n5563, \REG.mem_0_3 , 
        n5561, n15859, n15115, n13300, n13301, n15847, n15109, 
        n13298, n13297, n13264, n13265, n15841, n14551, n13259, 
        n13258, n13375, n13376, n15103, n14554, n13370, n13369, 
        n15829, n13861, n13862, n15097, n15823, n13118, n13117, 
        n15817, n15091, n15805, n15085, n13608, n13607, n13560, 
        n13559, n13776, n13775;
    
    SB_LUT4 i4722_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_18_22 ), .O(n6196));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4722_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4721_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_18_21 ), .O(n6195));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4721_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11126_3_lut (.I0(\REG.mem_0_9 ), .I1(\REG.mem_1_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13237));
    defparam i11126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11127_3_lut (.I0(\REG.mem_2_9 ), .I1(\REG.mem_3_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13238));
    defparam i11127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4720_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_18_20 ), .O(n6194));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4720_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14647_bdd_4_lut (.I0(n14647), .I1(n13064), .I2(n13063), .I3(rd_addr_r[2]), 
            .O(n14650));
    defparam n14647_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4719_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_18_19 ), .O(n6193));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4719_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4718_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_18_18 ), .O(n6192));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4718_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4717_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_18_17 ), .O(n6191));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4717_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11133_3_lut (.I0(\REG.mem_6_9 ), .I1(\REG.mem_7_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13244));
    defparam i11133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11132_3_lut (.I0(\REG.mem_4_9 ), .I1(\REG.mem_5_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13243));
    defparam i11132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4716_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_18_16 ), .O(n6190));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4716_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11159_3_lut (.I0(\REG.mem_24_9 ), .I1(\REG.mem_25_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13270));
    defparam i11159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13471 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_25 ), 
            .I2(\REG.mem_19_25 ), .I3(rd_addr_r[1]), .O(n15793));
    defparam rd_addr_r_0__bdd_4_lut_13471.LUT_INIT = 16'he4aa;
    SB_LUT4 n14515_bdd_4_lut (.I0(n14515), .I1(\REG.mem_1_31 ), .I2(\REG.mem_0_31 ), 
            .I3(rd_addr_r[1]), .O(n14518));
    defparam n14515_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15073_bdd_4_lut (.I0(n15073), .I1(\REG.mem_9_5 ), .I2(\REG.mem_8_5 ), 
            .I3(rd_addr_r[1]), .O(n14016));
    defparam n15073_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11160_3_lut (.I0(\REG.mem_26_9 ), .I1(\REG.mem_27_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13271));
    defparam i11160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i6_1_lut (.I0(rd_grey_sync_r[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n1[5]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n15793_bdd_4_lut (.I0(n15793), .I1(\REG.mem_17_25 ), .I2(\REG.mem_16_25 ), 
            .I3(rd_addr_r[1]), .O(n13794));
    defparam n15793_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4715_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_18_15 ), .O(n6189));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4715_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13461 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_16 ), 
            .I2(\REG.mem_7_16 ), .I3(rd_addr_r[1]), .O(n15787));
    defparam rd_addr_r_0__bdd_4_lut_13461.LUT_INIT = 16'he4aa;
    SB_LUT4 i11477_3_lut (.I0(\REG.mem_0_7 ), .I1(\REG.mem_1_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13588));
    defparam i11477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11478_3_lut (.I0(\REG.mem_2_7 ), .I1(\REG.mem_3_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13589));
    defparam i11478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4714_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_18_14 ), .O(n6188));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4714_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i25_2_lut_3_lut (.I0(n8_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n25_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i25_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i11130_3_lut (.I0(\REG.mem_6_7 ), .I1(\REG.mem_7_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13241));
    defparam i11130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11129_3_lut (.I0(\REG.mem_4_7 ), .I1(\REG.mem_5_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13240));
    defparam i11129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11166_3_lut (.I0(\REG.mem_30_9 ), .I1(\REG.mem_31_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13277));
    defparam i11166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12523 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_23 ), 
            .I2(\REG.mem_11_23 ), .I3(rd_addr_r[1]), .O(n14641));
    defparam rd_addr_r_0__bdd_4_lut_12523.LUT_INIT = 16'he4aa;
    SB_LUT4 i4713_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_18_13 ), .O(n6187));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4713_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15787_bdd_4_lut (.I0(n15787), .I1(\REG.mem_5_16 ), .I2(\REG.mem_4_16 ), 
            .I3(rd_addr_r[1]), .O(n13812));
    defparam n15787_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11165_3_lut (.I0(\REG.mem_28_9 ), .I1(\REG.mem_29_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13276));
    defparam i11165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12882 (.I0(rd_addr_r[1]), .I1(n14194), 
            .I2(n14195), .I3(rd_addr_r[2]), .O(n15067));
    defparam rd_addr_r_1__bdd_4_lut_12882.LUT_INIT = 16'he4aa;
    SB_LUT4 i4712_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_18_12 ), .O(n6186));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4712_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11162_3_lut (.I0(\REG.mem_16_7 ), .I1(\REG.mem_17_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13273));
    defparam i11162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11163_3_lut (.I0(\REG.mem_18_7 ), .I1(\REG.mem_19_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13274));
    defparam i11163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11787_3_lut (.I0(\REG.mem_22_7 ), .I1(\REG.mem_23_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13898));
    defparam i11787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11786_3_lut (.I0(\REG.mem_20_7 ), .I1(\REG.mem_21_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13897));
    defparam i11786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n15067_bdd_4_lut (.I0(n15067), .I1(n14189), .I2(n14188), .I3(rd_addr_r[2]), 
            .O(n13157));
    defparam n15067_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14641_bdd_4_lut (.I0(n14641), .I1(\REG.mem_9_23 ), .I2(\REG.mem_8_23 ), 
            .I3(rd_addr_r[1]), .O(n14644));
    defparam n14641_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4711_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_18_11 ), .O(n6185));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4711_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i56_2_lut_3_lut_4_lut (.I0(n8_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n7));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i56_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i57_2_lut_3_lut_4_lut (.I0(n8_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n23));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i57_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_DFF i356_357 (.Q(\REG.mem_3_10 ), .C(FIFO_CLK_c), .D(n5704));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_13051 (.I0(rd_addr_r[2]), .I1(n13929), 
            .I2(n13938), .I3(rd_addr_r[3]), .O(n15061));
    defparam rd_addr_r_2__bdd_4_lut_13051.LUT_INIT = 16'he4aa;
    SB_LUT4 i4710_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_18_10 ), .O(n6184));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4710_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15061_bdd_4_lut (.I0(n15061), .I1(n13911), .I2(n13890), .I3(rd_addr_r[3]), 
            .O(n15064));
    defparam n15061_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR \afull_flag_impl.af_flag_ext_r_111  (.Q(DEBUG_1_c), .C(FIFO_CLK_c), 
            .D(\afull_flag_impl.af_flag_nxt_w ), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(410[29] 422[32])
    SB_LUT4 EnabledDecoder_2_i12_2_lut_3_lut_4_lut (.I0(wr_fifo_en_w), .I1(\wr_addr_r[0] ), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[1]), .O(n12_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i12_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i4709_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_18_9 ), .O(n6183));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4709_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i13_2_lut_3_lut_4_lut (.I0(wr_fifo_en_w), .I1(\wr_addr_r[0] ), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[1]), .O(n13_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i13_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i4708_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_18_8 ), .O(n6182));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4708_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i353_354 (.Q(\REG.mem_3_9 ), .C(FIFO_CLK_c), .D(n5703));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5083_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_29_31 ), .O(n6557));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5083_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4707_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_18_7 ), .O(n6181));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4707_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5082_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_29_30 ), .O(n6556));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5082_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13456 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_29 ), 
            .I2(\REG.mem_23_29 ), .I3(rd_addr_r[1]), .O(n15775));
    defparam rd_addr_r_0__bdd_4_lut_13456.LUT_INIT = 16'he4aa;
    SB_LUT4 i4706_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_18_6 ), .O(n6180));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4706_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12857 (.I0(rd_addr_r[1]), .I1(n13366), 
            .I2(n13367), .I3(rd_addr_r[2]), .O(n15055));
    defparam rd_addr_r_1__bdd_4_lut_12857.LUT_INIT = 16'he4aa;
    SB_LUT4 n15775_bdd_4_lut (.I0(n15775), .I1(\REG.mem_21_29 ), .I2(\REG.mem_20_29 ), 
            .I3(rd_addr_r[1]), .O(n15778));
    defparam n15775_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5081_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_29_29 ), .O(n6555));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5081_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i350_351 (.Q(\REG.mem_3_8 ), .C(FIFO_CLK_c), .D(n5702));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4705_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_18_5 ), .O(n6179));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4705_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4704_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_18_4 ), .O(n6178));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4704_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15055_bdd_4_lut (.I0(n15055), .I1(n13361), .I2(n13360), .I3(rd_addr_r[2]), 
            .O(n13483));
    defparam n15055_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13446 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_11 ), 
            .I2(\REG.mem_15_11 ), .I3(rd_addr_r[1]), .O(n15769));
    defparam rd_addr_r_0__bdd_4_lut_13446.LUT_INIT = 16'he4aa;
    SB_DFFE \REG.out_raw_i0_i1  (.Q(DEBUG_5_c_0), .C(SLM_CLK_c), .E(rd_fifo_en_w), 
            .D(rd_data_o_31__N_598[0]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_LUT4 i5080_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_29_28 ), .O(n6554));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5080_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12862 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_21 ), 
            .I2(\REG.mem_27_21 ), .I3(rd_addr_r[1]), .O(n15049));
    defparam rd_addr_r_0__bdd_4_lut_12862.LUT_INIT = 16'he4aa;
    SB_LUT4 i5079_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_29_27 ), .O(n6553));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5079_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15769_bdd_4_lut (.I0(n15769), .I1(\REG.mem_13_11 ), .I2(\REG.mem_12_11 ), 
            .I3(rd_addr_r[1]), .O(n15772));
    defparam n15769_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13441 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_25 ), 
            .I2(\REG.mem_27_25 ), .I3(rd_addr_r[1]), .O(n15763));
    defparam rd_addr_r_0__bdd_4_lut_13441.LUT_INIT = 16'he4aa;
    SB_LUT4 i4703_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_18_3 ), .O(n6177));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4703_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15763_bdd_4_lut (.I0(n15763), .I1(\REG.mem_25_25 ), .I2(\REG.mem_24_25 ), 
            .I3(rd_addr_r[1]), .O(n13827));
    defparam n15763_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15049_bdd_4_lut (.I0(n15049), .I1(\REG.mem_25_21 ), .I2(\REG.mem_24_21 ), 
            .I3(rd_addr_r[1]), .O(n15052));
    defparam n15049_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11177_3_lut (.I0(\REG.mem_0_10 ), .I1(\REG.mem_1_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13288));
    defparam i11177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11178_3_lut (.I0(\REG.mem_2_10 ), .I1(\REG.mem_3_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13289));
    defparam i11178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4702_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_18_2 ), .O(n6176));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4702_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4701_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_18_1 ), .O(n6175));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4701_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5078_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_29_26 ), .O(n6552));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5078_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4700_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_18_0 ), .O(n6174));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4700_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11184_3_lut (.I0(\REG.mem_6_10 ), .I1(\REG.mem_7_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13295));
    defparam i11184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11183_3_lut (.I0(\REG.mem_4_10 ), .I1(\REG.mem_5_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13294));
    defparam i11183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12842 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_26 ), 
            .I2(\REG.mem_3_26 ), .I3(rd_addr_r[1]), .O(n15043));
    defparam rd_addr_r_0__bdd_4_lut_12842.LUT_INIT = 16'he4aa;
    SB_LUT4 n15043_bdd_4_lut (.I0(n15043), .I1(\REG.mem_1_26 ), .I2(\REG.mem_0_26 ), 
            .I3(rd_addr_r[1]), .O(n15046));
    defparam n15043_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13436 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_16 ), 
            .I2(\REG.mem_15_16 ), .I3(rd_addr_r[1]), .O(n15757));
    defparam rd_addr_r_0__bdd_4_lut_13436.LUT_INIT = 16'he4aa;
    SB_LUT4 i5077_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_29_25 ), .O(n6551));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5077_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12852 (.I0(rd_addr_r[2]), .I1(n13944), 
            .I2(n13956), .I3(rd_addr_r[3]), .O(n15037));
    defparam rd_addr_r_2__bdd_4_lut_12852.LUT_INIT = 16'he4aa;
    SB_LUT4 n15037_bdd_4_lut (.I0(n15037), .I1(n13935), .I2(n13923), .I3(rd_addr_r[3]), 
            .O(n15040));
    defparam n15037_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15757_bdd_4_lut (.I0(n15757), .I1(\REG.mem_13_16 ), .I2(\REG.mem_12_16 ), 
            .I3(rd_addr_r[1]), .O(n13830));
    defparam n15757_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12837 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_5 ), 
            .I2(\REG.mem_15_5 ), .I3(rd_addr_r[1]), .O(n15031));
    defparam rd_addr_r_0__bdd_4_lut_12837.LUT_INIT = 16'he4aa;
    SB_LUT4 n15031_bdd_4_lut (.I0(n15031), .I1(\REG.mem_13_5 ), .I2(\REG.mem_12_5 ), 
            .I3(rd_addr_r[1]), .O(n14025));
    defparam n15031_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13501 (.I0(rd_addr_r[1]), .I1(n13309), 
            .I2(n13310), .I3(rd_addr_r[2]), .O(n15751));
    defparam rd_addr_r_1__bdd_4_lut_13501.LUT_INIT = 16'he4aa;
    SB_LUT4 n15751_bdd_4_lut (.I0(n15751), .I1(n13292), .I2(n13291), .I3(rd_addr_r[2]), 
            .O(n13837));
    defparam n15751_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i347_348 (.Q(\REG.mem_3_7 ), .C(FIFO_CLK_c), .D(n5701));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12832 (.I0(rd_addr_r[2]), .I1(n13986), 
            .I2(n13995), .I3(rd_addr_r[3]), .O(n15025));
    defparam rd_addr_r_2__bdd_4_lut_12832.LUT_INIT = 16'he4aa;
    SB_DFF i344_345 (.Q(\REG.mem_3_6 ), .C(FIFO_CLK_c), .D(n5700));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n15025_bdd_4_lut (.I0(n15025), .I1(n13971), .I2(n13953), .I3(rd_addr_r[3]), 
            .O(n15028));
    defparam n15025_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i47_2_lut_3_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n28));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i47_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i46_2_lut_3_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n12));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i46_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13431 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_29 ), 
            .I2(\REG.mem_15_29 ), .I3(rd_addr_r[1]), .O(n15745));
    defparam rd_addr_r_0__bdd_4_lut_13431.LUT_INIT = 16'he4aa;
    SB_LUT4 i5076_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_29_24 ), .O(n6550));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5076_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5075_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_29_23 ), .O(n6549));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5075_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15745_bdd_4_lut (.I0(n15745), .I1(\REG.mem_13_29 ), .I2(\REG.mem_12_29 ), 
            .I3(rd_addr_r[1]), .O(n15748));
    defparam n15745_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i341_342 (.Q(\REG.mem_3_5 ), .C(FIFO_CLK_c), .D(n5699));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFSR rd_grey_sync_r__i0 (.Q(rd_grey_sync_r[0]), .C(SLM_CLK_c), .D(rd_grey_w[0]), 
            .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12847 (.I0(rd_addr_r[1]), .I1(n13114), 
            .I2(n13115), .I3(rd_addr_r[2]), .O(n15019));
    defparam rd_addr_r_1__bdd_4_lut_12847.LUT_INIT = 16'he4aa;
    SB_DFFSS empty_ext_r_114 (.Q(dc32_fifo_empty), .C(SLM_CLK_c), .D(empty_nxt_c_N_636), 
            .S(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFFSR wr_grey_sync_r__i0 (.Q(\wr_grey_sync_r[0] ), .C(FIFO_CLK_c), 
            .D(wr_grey_w[0]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFF i338_339 (.Q(\REG.mem_3_4 ), .C(FIFO_CLK_c), .D(n5698));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFS \aempty_flag_impl.ae_flag_ext_r_120  (.Q(dc32_fifo_almost_empty), 
            .C(SLM_CLK_c), .D(\aempty_flag_impl.ae_flag_nxt_w ), .S(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(669[37] 672[40])
    SB_LUT4 i5074_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_29_22 ), .O(n6548));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5074_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12405 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_31 ), 
            .I2(\REG.mem_3_31 ), .I3(rd_addr_r[1]), .O(n14515));
    defparam rd_addr_r_0__bdd_4_lut_12405.LUT_INIT = 16'he4aa;
    SB_LUT4 i5073_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_29_21 ), .O(n6547));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5073_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5072_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_29_20 ), .O(n6546));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5072_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15019_bdd_4_lut (.I0(n15019), .I1(n13085), .I2(n13084), .I3(rd_addr_r[2]), 
            .O(n15022));
    defparam n15019_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i39_2_lut_3_lut (.I0(n15), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n32));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i39_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i38_2_lut_3_lut (.I0(n15), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n16));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i38_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i5071_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_29_19 ), .O(n6545));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5071_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13426 (.I0(rd_addr_r[1]), .I1(n13060), 
            .I2(n13061), .I3(rd_addr_r[2]), .O(n15721));
    defparam rd_addr_r_1__bdd_4_lut_13426.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12916 (.I0(rd_addr_r[3]), .I1(n14998), 
            .I2(n13436), .I3(rd_addr_r[4]), .O(n15013));
    defparam rd_addr_r_3__bdd_4_lut_12916.LUT_INIT = 16'he4aa;
    SB_LUT4 n15721_bdd_4_lut (.I0(n15721), .I1(n13322), .I2(n13321), .I3(rd_addr_r[2]), 
            .O(n13838));
    defparam n15721_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_13551 (.I0(rd_addr_r[3]), .I1(n13729), 
            .I2(n13730), .I3(rd_addr_r[4]), .O(n15715));
    defparam rd_addr_r_3__bdd_4_lut_13551.LUT_INIT = 16'he4aa;
    SB_LUT4 n15715_bdd_4_lut (.I0(n15715), .I1(n13694), .I2(n15496), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[29]));
    defparam n15715_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15013_bdd_4_lut (.I0(n15013), .I1(n13433), .I2(n14992), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[27]));
    defparam n15013_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13401 (.I0(rd_addr_r[1]), .I1(n13357), 
            .I2(n13358), .I3(rd_addr_r[2]), .O(n15709));
    defparam rd_addr_r_1__bdd_4_lut_13401.LUT_INIT = 16'he4aa;
    SB_LUT4 i5070_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_29_18 ), .O(n6544));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5070_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12817 (.I0(rd_addr_r[1]), .I1(n13402), 
            .I2(n13403), .I3(rd_addr_r[2]), .O(n15007));
    defparam rd_addr_r_1__bdd_4_lut_12817.LUT_INIT = 16'he4aa;
    SB_LUT4 n15007_bdd_4_lut (.I0(n15007), .I1(n13397), .I2(n13396), .I3(rd_addr_r[2]), 
            .O(n13444));
    defparam n15007_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5069_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_29_17 ), .O(n6543));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5069_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5068_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_29_16 ), .O(n6542));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5068_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5067_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_29_15 ), .O(n6541));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5067_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5066_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_29_14 ), .O(n6540));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5066_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5065_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_29_13 ), .O(n6539));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5065_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5064_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_29_12 ), .O(n6538));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5064_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12807 (.I0(rd_addr_r[1]), .I1(n13738), 
            .I2(n13739), .I3(rd_addr_r[2]), .O(n14995));
    defparam rd_addr_r_1__bdd_4_lut_12807.LUT_INIT = 16'he4aa;
    SB_DFF i335_336 (.Q(\REG.mem_3_3 ), .C(FIFO_CLK_c), .D(n5697));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n15709_bdd_4_lut (.I0(n15709), .I1(n13349), .I2(n13348), .I3(rd_addr_r[2]), 
            .O(n13379));
    defparam n15709_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14995_bdd_4_lut (.I0(n14995), .I1(n14174), .I2(n14173), .I3(rd_addr_r[2]), 
            .O(n14998));
    defparam n14995_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5063_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_29_11 ), .O(n6537));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5063_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5062_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_29_10 ), .O(n6536));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5062_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5061_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_29_9 ), .O(n6535));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5061_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12797 (.I0(rd_addr_r[1]), .I1(n14122), 
            .I2(n14123), .I3(rd_addr_r[2]), .O(n14989));
    defparam rd_addr_r_1__bdd_4_lut_12797.LUT_INIT = 16'he4aa;
    SB_LUT4 i5060_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_29_8 ), .O(n6534));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5060_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13421 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_25 ), 
            .I2(\REG.mem_31_25 ), .I3(rd_addr_r[1]), .O(n15691));
    defparam rd_addr_r_0__bdd_4_lut_13421.LUT_INIT = 16'he4aa;
    SB_DFF i332_333 (.Q(\REG.mem_3_2 ), .C(FIFO_CLK_c), .D(n5696));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i11579_3_lut (.I0(n15046), .I1(n14566), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13690));
    defparam i11579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n15691_bdd_4_lut (.I0(n15691), .I1(\REG.mem_29_25 ), .I2(\REG.mem_28_25 ), 
            .I3(rd_addr_r[1]), .O(n13851));
    defparam n15691_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5059_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_29_7 ), .O(n6533));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5059_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14989_bdd_4_lut (.I0(n14989), .I1(n13769), .I2(n13768), .I3(rd_addr_r[2]), 
            .O(n14992));
    defparam n14989_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13391 (.I0(rd_addr_r[1]), .I1(n13372), 
            .I2(n13373), .I3(rd_addr_r[2]), .O(n15685));
    defparam rd_addr_r_1__bdd_4_lut_13391.LUT_INIT = 16'he4aa;
    SB_LUT4 i10947_3_lut (.I0(n15862), .I1(n15598), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13058));
    defparam i10947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11195_3_lut (.I0(\REG.mem_16_10 ), .I1(\REG.mem_17_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13306));
    defparam i11195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11196_3_lut (.I0(\REG.mem_18_10 ), .I1(\REG.mem_19_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13307));
    defparam i11196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11202_3_lut (.I0(\REG.mem_22_10 ), .I1(\REG.mem_23_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13313));
    defparam i11202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11201_3_lut (.I0(\REG.mem_20_10 ), .I1(\REG.mem_21_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13312));
    defparam i11201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_2_lut (.I0(n7_adj_1372), .I1(n8_adj_1373), .I2(GND_net), 
            .I3(GND_net), .O(n12209));
    defparam i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 wr_addr_r_5__I_0_inv_0_i6_1_lut (.I0(rp_sync2_r[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1394[5]));   // src/fifo_dc_32_lut_gen.v(212[47:78])
    defparam wr_addr_r_5__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5058_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_29_6 ), .O(n6532));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5058_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4230_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_3_10 ), .O(n5704));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4230_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4229_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_3_9 ), .O(n5703));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4229_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4228_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_3_8 ), .O(n5702));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4228_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11741_3_lut (.I0(n14902), .I1(n15640), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13852));
    defparam i11741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4227_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_3_7 ), .O(n5701));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4227_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15685_bdd_4_lut (.I0(n15685), .I1(n13364), .I2(n13363), .I3(rd_addr_r[2]), 
            .O(n13391));
    defparam n15685_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4226_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_3_6 ), .O(n5700));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4226_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11742_3_lut (.I0(n15202), .I1(n16180), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13853));
    defparam i11742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4225_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_3_5 ), .O(n5699));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4225_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12812 (.I0(rd_addr_r[3]), .I1(n13444), 
            .I2(n13445), .I3(rd_addr_r[4]), .O(n14977));
    defparam rd_addr_r_3__bdd_4_lut_12812.LUT_INIT = 16'he4aa;
    SB_LUT4 i5057_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_29_5 ), .O(n6531));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5057_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4224_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_3_4 ), .O(n5698));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4224_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4223_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_3_3 ), .O(n5697));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4223_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4222_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_3_2 ), .O(n5696));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4222_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5056_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_29_4 ), .O(n6530));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5056_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5055_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_29_3 ), .O(n6529));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5055_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5054_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_29_2 ), .O(n6528));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5054_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4221_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_3_1 ), .O(n5695));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4221_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5053_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_29_1 ), .O(n6527));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5053_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14977_bdd_4_lut (.I0(n14977), .I1(n13418), .I2(n14968), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[1]));
    defparam n14977_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4220_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_3_0 ), .O(n5694));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4220_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4251_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_3_31 ), .O(n5725));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4251_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4250_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_3_30 ), .O(n5724));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4250_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4249_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_3_29 ), .O(n5723));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4249_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i329_330 (.Q(\REG.mem_3_1 ), .C(FIFO_CLK_c), .D(n5695));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i326_327 (.Q(\REG.mem_3_0 ), .C(FIFO_CLK_c), .D(n5694));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5052_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_29_0 ), .O(n6526));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5052_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFSR full_ext_r_107 (.Q(dc32_fifo_full), .C(FIFO_CLK_c), .D(full_nxt_c_N_633), 
            .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 i4248_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_3_28 ), .O(n5722));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4248_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12822 (.I0(rd_addr_r[2]), .I1(n14704), 
            .I2(n14692), .I3(rd_addr_r[3]), .O(n14971));
    defparam rd_addr_r_2__bdd_4_lut_12822.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13376 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_28 ), 
            .I2(\REG.mem_11_28 ), .I3(rd_addr_r[1]), .O(n15673));
    defparam rd_addr_r_0__bdd_4_lut_13376.LUT_INIT = 16'he4aa;
    SB_LUT4 i4247_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_3_27 ), .O(n5721));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4247_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14971_bdd_4_lut (.I0(n14971), .I1(n14722), .I2(n14764), .I3(rd_addr_r[3]), 
            .O(n14974));
    defparam n14971_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4246_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_3_26 ), .O(n5720));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4246_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15673_bdd_4_lut (.I0(n15673), .I1(\REG.mem_9_28 ), .I2(\REG.mem_8_28 ), 
            .I3(rd_addr_r[1]), .O(n15676));
    defparam n15673_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4245_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_3_25 ), .O(n5719));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4245_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4244_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_3_24 ), .O(n5718));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4244_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4243_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_3_23 ), .O(n5717));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4243_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4242_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_3_22 ), .O(n5716));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4242_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4241_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_3_21 ), .O(n5715));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4241_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13361 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_1 ), 
            .I2(\REG.mem_15_1 ), .I3(rd_addr_r[1]), .O(n15667));
    defparam rd_addr_r_0__bdd_4_lut_13361.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12503 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_29 ), 
            .I2(\REG.mem_19_29 ), .I3(rd_addr_r[1]), .O(n14629));
    defparam rd_addr_r_0__bdd_4_lut_12503.LUT_INIT = 16'he4aa;
    SB_LUT4 n14629_bdd_4_lut (.I0(n14629), .I1(\REG.mem_17_29 ), .I2(\REG.mem_16_29 ), 
            .I3(rd_addr_r[1]), .O(n14632));
    defparam n14629_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i323_324 (.Q(\REG.mem_2_31 ), .C(FIFO_CLK_c), .D(n5693));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4240_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_3_20 ), .O(n5714));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4240_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i28_2_lut (.I0(n12_c), .I1(wr_addr_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n28_adj_1375));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4239_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_3_19 ), .O(n5713));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4239_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15667_bdd_4_lut (.I0(n15667), .I1(\REG.mem_13_1 ), .I2(\REG.mem_12_1 ), 
            .I3(rd_addr_r[1]), .O(n15670));
    defparam n15667_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12508 (.I0(rd_addr_r[1]), .I1(n13492), 
            .I2(n13493), .I3(rd_addr_r[2]), .O(n14623));
    defparam rd_addr_r_1__bdd_4_lut_12508.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12792 (.I0(rd_addr_r[1]), .I1(n13387), 
            .I2(n13388), .I3(rd_addr_r[2]), .O(n14965));
    defparam rd_addr_r_1__bdd_4_lut_12792.LUT_INIT = 16'he4aa;
    SB_LUT4 n14623_bdd_4_lut (.I0(n14623), .I1(n13481), .I2(n13480), .I3(rd_addr_r[2]), 
            .O(n14626));
    defparam n14623_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4238_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_3_18 ), .O(n5712));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4238_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4237_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_3_17 ), .O(n5711));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4237_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4236_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_3_16 ), .O(n5710));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4236_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4235_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_3_15 ), .O(n5709));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4235_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4234_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_3_14 ), .O(n5708));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4234_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4233_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_3_13 ), .O(n5707));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4233_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4232_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_3_12 ), .O(n5706));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4232_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_nxt_c_5__I_0_138_i3_2_lut_4_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1_w[2]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_5__N_573[3] ), .O(rd_grey_w[2]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_5__I_0_138_i3_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4231_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_3_11 ), .O(n5705));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4231_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_nxt_c_5__I_0_138_i2_2_lut_4_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1_w[2]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_5__N_573[1] ), .O(rd_grey_w[1]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_5__I_0_138_i2_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i5527_2_lut_4_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1_w[2]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n7001));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i5527_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 EnabledDecoder_2_i27_2_lut_3_lut (.I0(n10_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n27_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i27_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i58_2_lut_3_lut_4_lut (.I0(n10_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n6));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i58_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i59_2_lut_3_lut_4_lut (.I0(n10_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n22));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i59_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i11675_3_lut (.I0(\REG.mem_0_28 ), .I1(\REG.mem_1_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13786));
    defparam i11675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11676_3_lut (.I0(\REG.mem_2_28 ), .I1(\REG.mem_3_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13787));
    defparam i11676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11685_3_lut (.I0(\REG.mem_6_28 ), .I1(\REG.mem_7_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13796));
    defparam i11685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11684_3_lut (.I0(\REG.mem_4_28 ), .I1(\REG.mem_5_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13795));
    defparam i11684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11228_3_lut (.I0(\REG.mem_0_2 ), .I1(\REG.mem_1_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13339));
    defparam i11228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11229_3_lut (.I0(\REG.mem_2_2 ), .I1(\REG.mem_3_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13340));
    defparam i11229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11232_3_lut (.I0(\REG.mem_6_2 ), .I1(\REG.mem_7_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13343));
    defparam i11232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11231_3_lut (.I0(\REG.mem_4_2 ), .I1(\REG.mem_5_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13342));
    defparam i11231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10976_3_lut (.I0(\REG.mem_0_22 ), .I1(\REG.mem_1_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13087));
    defparam i10976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10977_3_lut (.I0(\REG.mem_2_22 ), .I1(\REG.mem_3_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13088));
    defparam i10977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11034_3_lut (.I0(\REG.mem_6_22 ), .I1(\REG.mem_7_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13145));
    defparam i11034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11033_3_lut (.I0(\REG.mem_4_22 ), .I1(\REG.mem_5_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13144));
    defparam i11033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11574_3_lut (.I0(n15520), .I1(n15406), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13685));
    defparam i11574_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11630_3_lut (.I0(n14878), .I1(n16132), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13741));
    defparam i11630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11240_3_lut (.I0(\REG.mem_16_22 ), .I1(\REG.mem_17_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13351));
    defparam i11240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11241_3_lut (.I0(\REG.mem_18_22 ), .I1(\REG.mem_19_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13352));
    defparam i11241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i14_2_lut_3_lut_4_lut (.I0(wr_fifo_en_w), .I1(\wr_addr_r[0] ), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[1]), .O(n14));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i14_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i11244_3_lut (.I0(\REG.mem_22_22 ), .I1(\REG.mem_23_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13355));
    defparam i11244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11243_3_lut (.I0(\REG.mem_20_22 ), .I1(\REG.mem_21_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13354));
    defparam i11243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i15_2_lut_3_lut_4_lut (.I0(wr_fifo_en_w), .I1(\wr_addr_r[0] ), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[1]), .O(n15));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i15_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 rd_addr_nxt_c_5__I_0_138_i5_2_lut_4_lut (.I0(rd_grey_sync_r[5]), 
            .I1(rd_addr_p1_w[5]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_5__N_573[4] ), 
            .O(rd_grey_w[4]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_5__I_0_138_i5_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i5525_2_lut_4_lut (.I0(rd_grey_sync_r[5]), .I1(rd_addr_p1_w[5]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n6999));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i5525_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 rd_addr_r_5__I_0_i4_3_lut (.I0(rd_addr_r[3]), .I1(rd_addr_p1_w[3]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_5__N_573[3] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_5__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12423 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_23 ), 
            .I2(\REG.mem_19_23 ), .I3(rd_addr_r[1]), .O(n14533));
    defparam rd_addr_r_0__bdd_4_lut_12423.LUT_INIT = 16'he4aa;
    SB_LUT4 n14965_bdd_4_lut (.I0(n14965), .I1(n13385), .I2(n13384), .I3(rd_addr_r[2]), 
            .O(n14968));
    defparam n14965_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14521_bdd_4_lut (.I0(n14521), .I1(\REG.mem_5_18 ), .I2(\REG.mem_4_18 ), 
            .I3(rd_addr_r[1]), .O(n14524));
    defparam n14521_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_5__I_0_i5_3_lut (.I0(rd_addr_r[4]), .I1(rd_addr_p1_w[4]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_5__N_573[4] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_5__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12493 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_4 ), 
            .I2(\REG.mem_7_4 ), .I3(rd_addr_r[1]), .O(n14617));
    defparam rd_addr_r_0__bdd_4_lut_12493.LUT_INIT = 16'he4aa;
    SB_LUT4 i4603_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_14_31 ), .O(n6077));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4603_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12414 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_18 ), 
            .I2(\REG.mem_7_18 ), .I3(rd_addr_r[1]), .O(n14521));
    defparam rd_addr_r_0__bdd_4_lut_12414.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13356 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_8 ), 
            .I2(\REG.mem_11_8 ), .I3(rd_addr_r[1]), .O(n15655));
    defparam rd_addr_r_0__bdd_4_lut_13356.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12782 (.I0(rd_addr_r[3]), .I1(n14956), 
            .I2(n13391), .I3(rd_addr_r[4]), .O(n14959));
    defparam rd_addr_r_3__bdd_4_lut_12782.LUT_INIT = 16'he4aa;
    SB_LUT4 n15655_bdd_4_lut (.I0(n15655), .I1(\REG.mem_9_8 ), .I2(\REG.mem_8_8 ), 
            .I3(rd_addr_r[1]), .O(n15658));
    defparam n15655_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14959_bdd_4_lut (.I0(n14959), .I1(n13382), .I2(n14944), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[22]));
    defparam n14959_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14617_bdd_4_lut (.I0(n14617), .I1(\REG.mem_5_4 ), .I2(\REG.mem_4_4 ), 
            .I3(rd_addr_r[1]), .O(n14620));
    defparam n14617_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13346 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_21 ), 
            .I2(\REG.mem_3_21 ), .I3(rd_addr_r[1]), .O(n15649));
    defparam rd_addr_r_0__bdd_4_lut_13346.LUT_INIT = 16'he4aa;
    SB_LUT4 n15649_bdd_4_lut (.I0(n15649), .I1(\REG.mem_1_21 ), .I2(\REG.mem_0_21 ), 
            .I3(rd_addr_r[1]), .O(n15652));
    defparam n15649_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF wp_sync2_r__i5 (.Q(wp_sync2_r[5]), .C(SLM_CLK_c), .D(n7013));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i4 (.Q(wp_sync2_r[4]), .C(SLM_CLK_c), .D(n7012));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i3 (.Q(wp_sync2_r[3]), .C(SLM_CLK_c), .D(n7011));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i2 (.Q(wp_sync2_r[2]), .C(SLM_CLK_c), .D(n7010));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i1 (.Q(wp_sync2_r[1]), .C(SLM_CLK_c), .D(n7009));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i5 (.Q(wp_sync1_r[5]), .C(SLM_CLK_c), .D(n7008));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i4 (.Q(wp_sync1_r[4]), .C(SLM_CLK_c), .D(n7007));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i3 (.Q(wp_sync1_r[3]), .C(SLM_CLK_c), .D(n7006));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i2 (.Q(wp_sync1_r[2]), .C(SLM_CLK_c), .D(n7005));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i1 (.Q(wp_sync1_r[1]), .C(SLM_CLK_c), .D(n7004));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF rd_addr_r__i4 (.Q(rd_addr_r[4]), .C(SLM_CLK_c), .D(n7003));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i3 (.Q(rd_addr_r[3]), .C(SLM_CLK_c), .D(n7002));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i2 (.Q(rd_addr_r[2]), .C(SLM_CLK_c), .D(n7001));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i1 (.Q(rd_addr_r[1]), .C(SLM_CLK_c), .D(n7000));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_grey_sync_r__i5 (.Q(rd_grey_sync_r[5]), .C(SLM_CLK_c), .D(n6999));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFF rp_sync2_r__i5 (.Q(rp_sync2_r[5]), .C(FIFO_CLK_c), .D(n6998));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i4 (.Q(rp_sync2_r[4]), .C(FIFO_CLK_c), .D(n6997));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i3 (.Q(rp_sync2_r[3]), .C(FIFO_CLK_c), .D(n6996));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i2 (.Q(rp_sync2_r[2]), .C(FIFO_CLK_c), .D(n6995));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i1 (.Q(rp_sync2_r[1]), .C(FIFO_CLK_c), .D(n6994));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i5 (.Q(rp_sync1_r[5]), .C(FIFO_CLK_c), .D(n6993));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i4 (.Q(rp_sync1_r[4]), .C(FIFO_CLK_c), .D(n6992));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i3 (.Q(rp_sync1_r[3]), .C(FIFO_CLK_c), .D(n6991));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i2 (.Q(rp_sync1_r[2]), .C(FIFO_CLK_c), .D(n6990));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i1 (.Q(rp_sync1_r[1]), .C(FIFO_CLK_c), .D(n6989));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13341 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_13 ), 
            .I2(\REG.mem_3_13 ), .I3(rd_addr_r[1]), .O(n15643));
    defparam rd_addr_r_0__bdd_4_lut_13341.LUT_INIT = 16'he4aa;
    SB_LUT4 n15643_bdd_4_lut (.I0(n15643), .I1(\REG.mem_1_13 ), .I2(\REG.mem_0_13 ), 
            .I3(rd_addr_r[1]), .O(n13869));
    defparam n15643_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF wr_addr_r__i1 (.Q(wr_addr_r[1]), .C(FIFO_CLK_c), .D(n6931));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i2 (.Q(wr_addr_r[2]), .C(FIFO_CLK_c), .D(n6930));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i3 (.Q(wr_addr_r[3]), .C(FIFO_CLK_c), .D(n6929));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i4 (.Q(wr_addr_r[4]), .C(FIFO_CLK_c), .D(n6928));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i5 (.Q(\wr_addr_r[5] ), .C(FIFO_CLK_c), .D(n6927));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13336 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_30 ), 
            .I2(\REG.mem_7_30 ), .I3(rd_addr_r[1]), .O(n15637));
    defparam rd_addr_r_0__bdd_4_lut_13336.LUT_INIT = 16'he4aa;
    SB_DFF i3107_3108 (.Q(\REG.mem_31_31 ), .C(FIFO_CLK_c), .D(n6621));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3104_3105 (.Q(\REG.mem_31_30 ), .C(FIFO_CLK_c), .D(n6620));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3101_3102 (.Q(\REG.mem_31_29 ), .C(FIFO_CLK_c), .D(n6619));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3098_3099 (.Q(\REG.mem_31_28 ), .C(FIFO_CLK_c), .D(n6618));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3095_3096 (.Q(\REG.mem_31_27 ), .C(FIFO_CLK_c), .D(n6617));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3092_3093 (.Q(\REG.mem_31_26 ), .C(FIFO_CLK_c), .D(n6616));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3089_3090 (.Q(\REG.mem_31_25 ), .C(FIFO_CLK_c), .D(n6615));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3086_3087 (.Q(\REG.mem_31_24 ), .C(FIFO_CLK_c), .D(n6614));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3083_3084 (.Q(\REG.mem_31_23 ), .C(FIFO_CLK_c), .D(n6613));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3080_3081 (.Q(\REG.mem_31_22 ), .C(FIFO_CLK_c), .D(n6612));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3077_3078 (.Q(\REG.mem_31_21 ), .C(FIFO_CLK_c), .D(n6611));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3074_3075 (.Q(\REG.mem_31_20 ), .C(FIFO_CLK_c), .D(n6610));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3071_3072 (.Q(\REG.mem_31_19 ), .C(FIFO_CLK_c), .D(n6609));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3068_3069 (.Q(\REG.mem_31_18 ), .C(FIFO_CLK_c), .D(n6608));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3065_3066 (.Q(\REG.mem_31_17 ), .C(FIFO_CLK_c), .D(n6607));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3062_3063 (.Q(\REG.mem_31_16 ), .C(FIFO_CLK_c), .D(n6606));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3059_3060 (.Q(\REG.mem_31_15 ), .C(FIFO_CLK_c), .D(n6605));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3056_3057 (.Q(\REG.mem_31_14 ), .C(FIFO_CLK_c), .D(n6604));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3053_3054 (.Q(\REG.mem_31_13 ), .C(FIFO_CLK_c), .D(n6603));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3050_3051 (.Q(\REG.mem_31_12 ), .C(FIFO_CLK_c), .D(n6602));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3047_3048 (.Q(\REG.mem_31_11 ), .C(FIFO_CLK_c), .D(n6601));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3044_3045 (.Q(\REG.mem_31_10 ), .C(FIFO_CLK_c), .D(n6600));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3041_3042 (.Q(\REG.mem_31_9 ), .C(FIFO_CLK_c), .D(n6599));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3038_3039 (.Q(\REG.mem_31_8 ), .C(FIFO_CLK_c), .D(n6598));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3035_3036 (.Q(\REG.mem_31_7 ), .C(FIFO_CLK_c), .D(n6597));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3032_3033 (.Q(\REG.mem_31_6 ), .C(FIFO_CLK_c), .D(n6596));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3029_3030 (.Q(\REG.mem_31_5 ), .C(FIFO_CLK_c), .D(n6595));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3026_3027 (.Q(\REG.mem_31_4 ), .C(FIFO_CLK_c), .D(n6594));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3023_3024 (.Q(\REG.mem_31_3 ), .C(FIFO_CLK_c), .D(n6593));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3020_3021 (.Q(\REG.mem_31_2 ), .C(FIFO_CLK_c), .D(n6592));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3017_3018 (.Q(\REG.mem_31_1 ), .C(FIFO_CLK_c), .D(n6591));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3014_3015 (.Q(\REG.mem_31_0 ), .C(FIFO_CLK_c), .D(n6590));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3011_3012 (.Q(\REG.mem_30_31 ), .C(FIFO_CLK_c), .D(n6589));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3008_3009 (.Q(\REG.mem_30_30 ), .C(FIFO_CLK_c), .D(n6588));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3005_3006 (.Q(\REG.mem_30_29 ), .C(FIFO_CLK_c), .D(n6587));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3002_3003 (.Q(\REG.mem_30_28 ), .C(FIFO_CLK_c), .D(n6586));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2999_3000 (.Q(\REG.mem_30_27 ), .C(FIFO_CLK_c), .D(n6585));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2996_2997 (.Q(\REG.mem_30_26 ), .C(FIFO_CLK_c), .D(n6584));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2993_2994 (.Q(\REG.mem_30_25 ), .C(FIFO_CLK_c), .D(n6583));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2990_2991 (.Q(\REG.mem_30_24 ), .C(FIFO_CLK_c), .D(n6582));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2987_2988 (.Q(\REG.mem_30_23 ), .C(FIFO_CLK_c), .D(n6581));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2984_2985 (.Q(\REG.mem_30_22 ), .C(FIFO_CLK_c), .D(n6580));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2981_2982 (.Q(\REG.mem_30_21 ), .C(FIFO_CLK_c), .D(n6579));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2978_2979 (.Q(\REG.mem_30_20 ), .C(FIFO_CLK_c), .D(n6578));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2975_2976 (.Q(\REG.mem_30_19 ), .C(FIFO_CLK_c), .D(n6577));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2972_2973 (.Q(\REG.mem_30_18 ), .C(FIFO_CLK_c), .D(n6576));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2969_2970 (.Q(\REG.mem_30_17 ), .C(FIFO_CLK_c), .D(n6575));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2966_2967 (.Q(\REG.mem_30_16 ), .C(FIFO_CLK_c), .D(n6574));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2963_2964 (.Q(\REG.mem_30_15 ), .C(FIFO_CLK_c), .D(n6573));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2960_2961 (.Q(\REG.mem_30_14 ), .C(FIFO_CLK_c), .D(n6572));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2957_2958 (.Q(\REG.mem_30_13 ), .C(FIFO_CLK_c), .D(n6571));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2954_2955 (.Q(\REG.mem_30_12 ), .C(FIFO_CLK_c), .D(n6570));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2951_2952 (.Q(\REG.mem_30_11 ), .C(FIFO_CLK_c), .D(n6569));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2948_2949 (.Q(\REG.mem_30_10 ), .C(FIFO_CLK_c), .D(n6568));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2945_2946 (.Q(\REG.mem_30_9 ), .C(FIFO_CLK_c), .D(n6567));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2942_2943 (.Q(\REG.mem_30_8 ), .C(FIFO_CLK_c), .D(n6566));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2939_2940 (.Q(\REG.mem_30_7 ), .C(FIFO_CLK_c), .D(n6565));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2936_2937 (.Q(\REG.mem_30_6 ), .C(FIFO_CLK_c), .D(n6564));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2933_2934 (.Q(\REG.mem_30_5 ), .C(FIFO_CLK_c), .D(n6563));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2930_2931 (.Q(\REG.mem_30_4 ), .C(FIFO_CLK_c), .D(n6562));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2927_2928 (.Q(\REG.mem_30_3 ), .C(FIFO_CLK_c), .D(n6561));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2924_2925 (.Q(\REG.mem_30_2 ), .C(FIFO_CLK_c), .D(n6560));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2921_2922 (.Q(\REG.mem_30_1 ), .C(FIFO_CLK_c), .D(n6559));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2918_2919 (.Q(\REG.mem_30_0 ), .C(FIFO_CLK_c), .D(n6558));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2915_2916 (.Q(\REG.mem_29_31 ), .C(FIFO_CLK_c), .D(n6557));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2912_2913 (.Q(\REG.mem_29_30 ), .C(FIFO_CLK_c), .D(n6556));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2909_2910 (.Q(\REG.mem_29_29 ), .C(FIFO_CLK_c), .D(n6555));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2906_2907 (.Q(\REG.mem_29_28 ), .C(FIFO_CLK_c), .D(n6554));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2903_2904 (.Q(\REG.mem_29_27 ), .C(FIFO_CLK_c), .D(n6553));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2900_2901 (.Q(\REG.mem_29_26 ), .C(FIFO_CLK_c), .D(n6552));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2897_2898 (.Q(\REG.mem_29_25 ), .C(FIFO_CLK_c), .D(n6551));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2894_2895 (.Q(\REG.mem_29_24 ), .C(FIFO_CLK_c), .D(n6550));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2891_2892 (.Q(\REG.mem_29_23 ), .C(FIFO_CLK_c), .D(n6549));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2888_2889 (.Q(\REG.mem_29_22 ), .C(FIFO_CLK_c), .D(n6548));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2885_2886 (.Q(\REG.mem_29_21 ), .C(FIFO_CLK_c), .D(n6547));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2882_2883 (.Q(\REG.mem_29_20 ), .C(FIFO_CLK_c), .D(n6546));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2879_2880 (.Q(\REG.mem_29_19 ), .C(FIFO_CLK_c), .D(n6545));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2876_2877 (.Q(\REG.mem_29_18 ), .C(FIFO_CLK_c), .D(n6544));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2873_2874 (.Q(\REG.mem_29_17 ), .C(FIFO_CLK_c), .D(n6543));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2870_2871 (.Q(\REG.mem_29_16 ), .C(FIFO_CLK_c), .D(n6542));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2867_2868 (.Q(\REG.mem_29_15 ), .C(FIFO_CLK_c), .D(n6541));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2864_2865 (.Q(\REG.mem_29_14 ), .C(FIFO_CLK_c), .D(n6540));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2861_2862 (.Q(\REG.mem_29_13 ), .C(FIFO_CLK_c), .D(n6539));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2858_2859 (.Q(\REG.mem_29_12 ), .C(FIFO_CLK_c), .D(n6538));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2855_2856 (.Q(\REG.mem_29_11 ), .C(FIFO_CLK_c), .D(n6537));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2852_2853 (.Q(\REG.mem_29_10 ), .C(FIFO_CLK_c), .D(n6536));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2849_2850 (.Q(\REG.mem_29_9 ), .C(FIFO_CLK_c), .D(n6535));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2846_2847 (.Q(\REG.mem_29_8 ), .C(FIFO_CLK_c), .D(n6534));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2843_2844 (.Q(\REG.mem_29_7 ), .C(FIFO_CLK_c), .D(n6533));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2840_2841 (.Q(\REG.mem_29_6 ), .C(FIFO_CLK_c), .D(n6532));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2837_2838 (.Q(\REG.mem_29_5 ), .C(FIFO_CLK_c), .D(n6531));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2834_2835 (.Q(\REG.mem_29_4 ), .C(FIFO_CLK_c), .D(n6530));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2831_2832 (.Q(\REG.mem_29_3 ), .C(FIFO_CLK_c), .D(n6529));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2828_2829 (.Q(\REG.mem_29_2 ), .C(FIFO_CLK_c), .D(n6528));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2825_2826 (.Q(\REG.mem_29_1 ), .C(FIFO_CLK_c), .D(n6527));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2822_2823 (.Q(\REG.mem_29_0 ), .C(FIFO_CLK_c), .D(n6526));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2819_2820 (.Q(\REG.mem_28_31 ), .C(FIFO_CLK_c), .D(n6525));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2816_2817 (.Q(\REG.mem_28_30 ), .C(FIFO_CLK_c), .D(n6524));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2813_2814 (.Q(\REG.mem_28_29 ), .C(FIFO_CLK_c), .D(n6523));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2810_2811 (.Q(\REG.mem_28_28 ), .C(FIFO_CLK_c), .D(n6522));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2807_2808 (.Q(\REG.mem_28_27 ), .C(FIFO_CLK_c), .D(n6521));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2804_2805 (.Q(\REG.mem_28_26 ), .C(FIFO_CLK_c), .D(n6520));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2801_2802 (.Q(\REG.mem_28_25 ), .C(FIFO_CLK_c), .D(n6519));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2798_2799 (.Q(\REG.mem_28_24 ), .C(FIFO_CLK_c), .D(n6518));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2795_2796 (.Q(\REG.mem_28_23 ), .C(FIFO_CLK_c), .D(n6517));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2792_2793 (.Q(\REG.mem_28_22 ), .C(FIFO_CLK_c), .D(n6516));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2789_2790 (.Q(\REG.mem_28_21 ), .C(FIFO_CLK_c), .D(n6515));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2786_2787 (.Q(\REG.mem_28_20 ), .C(FIFO_CLK_c), .D(n6514));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2783_2784 (.Q(\REG.mem_28_19 ), .C(FIFO_CLK_c), .D(n6513));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2780_2781 (.Q(\REG.mem_28_18 ), .C(FIFO_CLK_c), .D(n6512));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2777_2778 (.Q(\REG.mem_28_17 ), .C(FIFO_CLK_c), .D(n6511));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2774_2775 (.Q(\REG.mem_28_16 ), .C(FIFO_CLK_c), .D(n6510));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2771_2772 (.Q(\REG.mem_28_15 ), .C(FIFO_CLK_c), .D(n6509));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2768_2769 (.Q(\REG.mem_28_14 ), .C(FIFO_CLK_c), .D(n6508));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2765_2766 (.Q(\REG.mem_28_13 ), .C(FIFO_CLK_c), .D(n6507));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2762_2763 (.Q(\REG.mem_28_12 ), .C(FIFO_CLK_c), .D(n6506));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2759_2760 (.Q(\REG.mem_28_11 ), .C(FIFO_CLK_c), .D(n6505));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2756_2757 (.Q(\REG.mem_28_10 ), .C(FIFO_CLK_c), .D(n6504));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2753_2754 (.Q(\REG.mem_28_9 ), .C(FIFO_CLK_c), .D(n6503));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2750_2751 (.Q(\REG.mem_28_8 ), .C(FIFO_CLK_c), .D(n6502));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2747_2748 (.Q(\REG.mem_28_7 ), .C(FIFO_CLK_c), .D(n6501));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2744_2745 (.Q(\REG.mem_28_6 ), .C(FIFO_CLK_c), .D(n6500));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2741_2742 (.Q(\REG.mem_28_5 ), .C(FIFO_CLK_c), .D(n6499));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2738_2739 (.Q(\REG.mem_28_4 ), .C(FIFO_CLK_c), .D(n6498));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2735_2736 (.Q(\REG.mem_28_3 ), .C(FIFO_CLK_c), .D(n6497));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2732_2733 (.Q(\REG.mem_28_2 ), .C(FIFO_CLK_c), .D(n6496));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2729_2730 (.Q(\REG.mem_28_1 ), .C(FIFO_CLK_c), .D(n6495));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2726_2727 (.Q(\REG.mem_28_0 ), .C(FIFO_CLK_c), .D(n6494));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2723_2724 (.Q(\REG.mem_27_31 ), .C(FIFO_CLK_c), .D(n6493));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2720_2721 (.Q(\REG.mem_27_30 ), .C(FIFO_CLK_c), .D(n6492));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2717_2718 (.Q(\REG.mem_27_29 ), .C(FIFO_CLK_c), .D(n6491));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2714_2715 (.Q(\REG.mem_27_28 ), .C(FIFO_CLK_c), .D(n6490));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2711_2712 (.Q(\REG.mem_27_27 ), .C(FIFO_CLK_c), .D(n6489));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2708_2709 (.Q(\REG.mem_27_26 ), .C(FIFO_CLK_c), .D(n6488));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2705_2706 (.Q(\REG.mem_27_25 ), .C(FIFO_CLK_c), .D(n6487));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2702_2703 (.Q(\REG.mem_27_24 ), .C(FIFO_CLK_c), .D(n6486));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2699_2700 (.Q(\REG.mem_27_23 ), .C(FIFO_CLK_c), .D(n6485));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2696_2697 (.Q(\REG.mem_27_22 ), .C(FIFO_CLK_c), .D(n6484));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2693_2694 (.Q(\REG.mem_27_21 ), .C(FIFO_CLK_c), .D(n6483));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2690_2691 (.Q(\REG.mem_27_20 ), .C(FIFO_CLK_c), .D(n6482));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2687_2688 (.Q(\REG.mem_27_19 ), .C(FIFO_CLK_c), .D(n6481));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2684_2685 (.Q(\REG.mem_27_18 ), .C(FIFO_CLK_c), .D(n6480));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2681_2682 (.Q(\REG.mem_27_17 ), .C(FIFO_CLK_c), .D(n6479));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2678_2679 (.Q(\REG.mem_27_16 ), .C(FIFO_CLK_c), .D(n6478));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2675_2676 (.Q(\REG.mem_27_15 ), .C(FIFO_CLK_c), .D(n6477));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2672_2673 (.Q(\REG.mem_27_14 ), .C(FIFO_CLK_c), .D(n6476));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2669_2670 (.Q(\REG.mem_27_13 ), .C(FIFO_CLK_c), .D(n6475));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2666_2667 (.Q(\REG.mem_27_12 ), .C(FIFO_CLK_c), .D(n6474));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2663_2664 (.Q(\REG.mem_27_11 ), .C(FIFO_CLK_c), .D(n6473));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2660_2661 (.Q(\REG.mem_27_10 ), .C(FIFO_CLK_c), .D(n6472));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2657_2658 (.Q(\REG.mem_27_9 ), .C(FIFO_CLK_c), .D(n6471));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2654_2655 (.Q(\REG.mem_27_8 ), .C(FIFO_CLK_c), .D(n6470));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2651_2652 (.Q(\REG.mem_27_7 ), .C(FIFO_CLK_c), .D(n6469));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2648_2649 (.Q(\REG.mem_27_6 ), .C(FIFO_CLK_c), .D(n6468));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2645_2646 (.Q(\REG.mem_27_5 ), .C(FIFO_CLK_c), .D(n6467));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2642_2643 (.Q(\REG.mem_27_4 ), .C(FIFO_CLK_c), .D(n6466));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2639_2640 (.Q(\REG.mem_27_3 ), .C(FIFO_CLK_c), .D(n6465));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2636_2637 (.Q(\REG.mem_27_2 ), .C(FIFO_CLK_c), .D(n6464));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2633_2634 (.Q(\REG.mem_27_1 ), .C(FIFO_CLK_c), .D(n6463));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2630_2631 (.Q(\REG.mem_27_0 ), .C(FIFO_CLK_c), .D(n6462));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2627_2628 (.Q(\REG.mem_26_31 ), .C(FIFO_CLK_c), .D(n6461));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2624_2625 (.Q(\REG.mem_26_30 ), .C(FIFO_CLK_c), .D(n6460));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2621_2622 (.Q(\REG.mem_26_29 ), .C(FIFO_CLK_c), .D(n6459));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2618_2619 (.Q(\REG.mem_26_28 ), .C(FIFO_CLK_c), .D(n6458));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2615_2616 (.Q(\REG.mem_26_27 ), .C(FIFO_CLK_c), .D(n6457));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2612_2613 (.Q(\REG.mem_26_26 ), .C(FIFO_CLK_c), .D(n6456));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2609_2610 (.Q(\REG.mem_26_25 ), .C(FIFO_CLK_c), .D(n6455));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2606_2607 (.Q(\REG.mem_26_24 ), .C(FIFO_CLK_c), .D(n6454));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2603_2604 (.Q(\REG.mem_26_23 ), .C(FIFO_CLK_c), .D(n6453));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2600_2601 (.Q(\REG.mem_26_22 ), .C(FIFO_CLK_c), .D(n6452));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2597_2598 (.Q(\REG.mem_26_21 ), .C(FIFO_CLK_c), .D(n6451));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2594_2595 (.Q(\REG.mem_26_20 ), .C(FIFO_CLK_c), .D(n6450));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2591_2592 (.Q(\REG.mem_26_19 ), .C(FIFO_CLK_c), .D(n6449));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2588_2589 (.Q(\REG.mem_26_18 ), .C(FIFO_CLK_c), .D(n6448));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2585_2586 (.Q(\REG.mem_26_17 ), .C(FIFO_CLK_c), .D(n6447));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2582_2583 (.Q(\REG.mem_26_16 ), .C(FIFO_CLK_c), .D(n6446));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2579_2580 (.Q(\REG.mem_26_15 ), .C(FIFO_CLK_c), .D(n6445));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2576_2577 (.Q(\REG.mem_26_14 ), .C(FIFO_CLK_c), .D(n6444));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2573_2574 (.Q(\REG.mem_26_13 ), .C(FIFO_CLK_c), .D(n6443));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2570_2571 (.Q(\REG.mem_26_12 ), .C(FIFO_CLK_c), .D(n6442));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2567_2568 (.Q(\REG.mem_26_11 ), .C(FIFO_CLK_c), .D(n6441));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2564_2565 (.Q(\REG.mem_26_10 ), .C(FIFO_CLK_c), .D(n6440));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2561_2562 (.Q(\REG.mem_26_9 ), .C(FIFO_CLK_c), .D(n6439));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2558_2559 (.Q(\REG.mem_26_8 ), .C(FIFO_CLK_c), .D(n6438));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2555_2556 (.Q(\REG.mem_26_7 ), .C(FIFO_CLK_c), .D(n6437));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2552_2553 (.Q(\REG.mem_26_6 ), .C(FIFO_CLK_c), .D(n6436));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2549_2550 (.Q(\REG.mem_26_5 ), .C(FIFO_CLK_c), .D(n6435));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2546_2547 (.Q(\REG.mem_26_4 ), .C(FIFO_CLK_c), .D(n6434));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2543_2544 (.Q(\REG.mem_26_3 ), .C(FIFO_CLK_c), .D(n6433));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2540_2541 (.Q(\REG.mem_26_2 ), .C(FIFO_CLK_c), .D(n6432));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2537_2538 (.Q(\REG.mem_26_1 ), .C(FIFO_CLK_c), .D(n6431));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2534_2535 (.Q(\REG.mem_26_0 ), .C(FIFO_CLK_c), .D(n6430));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2531_2532 (.Q(\REG.mem_25_31 ), .C(FIFO_CLK_c), .D(n6429));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2528_2529 (.Q(\REG.mem_25_30 ), .C(FIFO_CLK_c), .D(n6428));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2525_2526 (.Q(\REG.mem_25_29 ), .C(FIFO_CLK_c), .D(n6427));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2522_2523 (.Q(\REG.mem_25_28 ), .C(FIFO_CLK_c), .D(n6426));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2519_2520 (.Q(\REG.mem_25_27 ), .C(FIFO_CLK_c), .D(n6425));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2516_2517 (.Q(\REG.mem_25_26 ), .C(FIFO_CLK_c), .D(n6424));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2513_2514 (.Q(\REG.mem_25_25 ), .C(FIFO_CLK_c), .D(n6423));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2510_2511 (.Q(\REG.mem_25_24 ), .C(FIFO_CLK_c), .D(n6422));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2507_2508 (.Q(\REG.mem_25_23 ), .C(FIFO_CLK_c), .D(n6421));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2504_2505 (.Q(\REG.mem_25_22 ), .C(FIFO_CLK_c), .D(n6420));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2501_2502 (.Q(\REG.mem_25_21 ), .C(FIFO_CLK_c), .D(n6419));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2498_2499 (.Q(\REG.mem_25_20 ), .C(FIFO_CLK_c), .D(n6418));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2495_2496 (.Q(\REG.mem_25_19 ), .C(FIFO_CLK_c), .D(n6417));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2492_2493 (.Q(\REG.mem_25_18 ), .C(FIFO_CLK_c), .D(n6416));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2489_2490 (.Q(\REG.mem_25_17 ), .C(FIFO_CLK_c), .D(n6415));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2486_2487 (.Q(\REG.mem_25_16 ), .C(FIFO_CLK_c), .D(n6414));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2483_2484 (.Q(\REG.mem_25_15 ), .C(FIFO_CLK_c), .D(n6413));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2480_2481 (.Q(\REG.mem_25_14 ), .C(FIFO_CLK_c), .D(n6412));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2477_2478 (.Q(\REG.mem_25_13 ), .C(FIFO_CLK_c), .D(n6411));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2474_2475 (.Q(\REG.mem_25_12 ), .C(FIFO_CLK_c), .D(n6410));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2471_2472 (.Q(\REG.mem_25_11 ), .C(FIFO_CLK_c), .D(n6409));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2468_2469 (.Q(\REG.mem_25_10 ), .C(FIFO_CLK_c), .D(n6408));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2465_2466 (.Q(\REG.mem_25_9 ), .C(FIFO_CLK_c), .D(n6407));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2462_2463 (.Q(\REG.mem_25_8 ), .C(FIFO_CLK_c), .D(n6406));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2459_2460 (.Q(\REG.mem_25_7 ), .C(FIFO_CLK_c), .D(n6405));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2456_2457 (.Q(\REG.mem_25_6 ), .C(FIFO_CLK_c), .D(n6404));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2453_2454 (.Q(\REG.mem_25_5 ), .C(FIFO_CLK_c), .D(n6403));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2450_2451 (.Q(\REG.mem_25_4 ), .C(FIFO_CLK_c), .D(n6402));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2447_2448 (.Q(\REG.mem_25_3 ), .C(FIFO_CLK_c), .D(n6401));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2444_2445 (.Q(\REG.mem_25_2 ), .C(FIFO_CLK_c), .D(n6400));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2441_2442 (.Q(\REG.mem_25_1 ), .C(FIFO_CLK_c), .D(n6399));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2438_2439 (.Q(\REG.mem_25_0 ), .C(FIFO_CLK_c), .D(n6398));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2435_2436 (.Q(\REG.mem_24_31 ), .C(FIFO_CLK_c), .D(n6397));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2432_2433 (.Q(\REG.mem_24_30 ), .C(FIFO_CLK_c), .D(n6396));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2429_2430 (.Q(\REG.mem_24_29 ), .C(FIFO_CLK_c), .D(n6395));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2426_2427 (.Q(\REG.mem_24_28 ), .C(FIFO_CLK_c), .D(n6394));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2423_2424 (.Q(\REG.mem_24_27 ), .C(FIFO_CLK_c), .D(n6393));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2420_2421 (.Q(\REG.mem_24_26 ), .C(FIFO_CLK_c), .D(n6392));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2417_2418 (.Q(\REG.mem_24_25 ), .C(FIFO_CLK_c), .D(n6391));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2414_2415 (.Q(\REG.mem_24_24 ), .C(FIFO_CLK_c), .D(n6390));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2411_2412 (.Q(\REG.mem_24_23 ), .C(FIFO_CLK_c), .D(n6389));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2408_2409 (.Q(\REG.mem_24_22 ), .C(FIFO_CLK_c), .D(n6388));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2405_2406 (.Q(\REG.mem_24_21 ), .C(FIFO_CLK_c), .D(n6387));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2402_2403 (.Q(\REG.mem_24_20 ), .C(FIFO_CLK_c), .D(n6386));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2399_2400 (.Q(\REG.mem_24_19 ), .C(FIFO_CLK_c), .D(n6385));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2396_2397 (.Q(\REG.mem_24_18 ), .C(FIFO_CLK_c), .D(n6384));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2393_2394 (.Q(\REG.mem_24_17 ), .C(FIFO_CLK_c), .D(n6383));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2390_2391 (.Q(\REG.mem_24_16 ), .C(FIFO_CLK_c), .D(n6382));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2387_2388 (.Q(\REG.mem_24_15 ), .C(FIFO_CLK_c), .D(n6381));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2384_2385 (.Q(\REG.mem_24_14 ), .C(FIFO_CLK_c), .D(n6380));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2381_2382 (.Q(\REG.mem_24_13 ), .C(FIFO_CLK_c), .D(n6379));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2378_2379 (.Q(\REG.mem_24_12 ), .C(FIFO_CLK_c), .D(n6378));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2375_2376 (.Q(\REG.mem_24_11 ), .C(FIFO_CLK_c), .D(n6377));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2372_2373 (.Q(\REG.mem_24_10 ), .C(FIFO_CLK_c), .D(n6376));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2369_2370 (.Q(\REG.mem_24_9 ), .C(FIFO_CLK_c), .D(n6375));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2366_2367 (.Q(\REG.mem_24_8 ), .C(FIFO_CLK_c), .D(n6374));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2363_2364 (.Q(\REG.mem_24_7 ), .C(FIFO_CLK_c), .D(n6373));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2360_2361 (.Q(\REG.mem_24_6 ), .C(FIFO_CLK_c), .D(n6372));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2357_2358 (.Q(\REG.mem_24_5 ), .C(FIFO_CLK_c), .D(n6371));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2354_2355 (.Q(\REG.mem_24_4 ), .C(FIFO_CLK_c), .D(n6370));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2351_2352 (.Q(\REG.mem_24_3 ), .C(FIFO_CLK_c), .D(n6369));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2348_2349 (.Q(\REG.mem_24_2 ), .C(FIFO_CLK_c), .D(n6368));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2345_2346 (.Q(\REG.mem_24_1 ), .C(FIFO_CLK_c), .D(n6367));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2342_2343 (.Q(\REG.mem_24_0 ), .C(FIFO_CLK_c), .D(n6366));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2339_2340 (.Q(\REG.mem_23_31 ), .C(FIFO_CLK_c), .D(n6365));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2336_2337 (.Q(\REG.mem_23_30 ), .C(FIFO_CLK_c), .D(n6364));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2333_2334 (.Q(\REG.mem_23_29 ), .C(FIFO_CLK_c), .D(n6363));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2330_2331 (.Q(\REG.mem_23_28 ), .C(FIFO_CLK_c), .D(n6362));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2327_2328 (.Q(\REG.mem_23_27 ), .C(FIFO_CLK_c), .D(n6361));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2324_2325 (.Q(\REG.mem_23_26 ), .C(FIFO_CLK_c), .D(n6360));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2321_2322 (.Q(\REG.mem_23_25 ), .C(FIFO_CLK_c), .D(n6359));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2318_2319 (.Q(\REG.mem_23_24 ), .C(FIFO_CLK_c), .D(n6358));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2315_2316 (.Q(\REG.mem_23_23 ), .C(FIFO_CLK_c), .D(n6357));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2312_2313 (.Q(\REG.mem_23_22 ), .C(FIFO_CLK_c), .D(n6356));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2309_2310 (.Q(\REG.mem_23_21 ), .C(FIFO_CLK_c), .D(n6355));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2306_2307 (.Q(\REG.mem_23_20 ), .C(FIFO_CLK_c), .D(n6354));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2303_2304 (.Q(\REG.mem_23_19 ), .C(FIFO_CLK_c), .D(n6353));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2300_2301 (.Q(\REG.mem_23_18 ), .C(FIFO_CLK_c), .D(n6352));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2297_2298 (.Q(\REG.mem_23_17 ), .C(FIFO_CLK_c), .D(n6351));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2294_2295 (.Q(\REG.mem_23_16 ), .C(FIFO_CLK_c), .D(n6350));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2291_2292 (.Q(\REG.mem_23_15 ), .C(FIFO_CLK_c), .D(n6349));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2288_2289 (.Q(\REG.mem_23_14 ), .C(FIFO_CLK_c), .D(n6348));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2285_2286 (.Q(\REG.mem_23_13 ), .C(FIFO_CLK_c), .D(n6347));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2282_2283 (.Q(\REG.mem_23_12 ), .C(FIFO_CLK_c), .D(n6346));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2279_2280 (.Q(\REG.mem_23_11 ), .C(FIFO_CLK_c), .D(n6345));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2276_2277 (.Q(\REG.mem_23_10 ), .C(FIFO_CLK_c), .D(n6344));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2273_2274 (.Q(\REG.mem_23_9 ), .C(FIFO_CLK_c), .D(n6343));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2270_2271 (.Q(\REG.mem_23_8 ), .C(FIFO_CLK_c), .D(n6342));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2267_2268 (.Q(\REG.mem_23_7 ), .C(FIFO_CLK_c), .D(n6341));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2264_2265 (.Q(\REG.mem_23_6 ), .C(FIFO_CLK_c), .D(n6340));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2261_2262 (.Q(\REG.mem_23_5 ), .C(FIFO_CLK_c), .D(n6339));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2258_2259 (.Q(\REG.mem_23_4 ), .C(FIFO_CLK_c), .D(n6338));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2255_2256 (.Q(\REG.mem_23_3 ), .C(FIFO_CLK_c), .D(n6337));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2252_2253 (.Q(\REG.mem_23_2 ), .C(FIFO_CLK_c), .D(n6336));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2249_2250 (.Q(\REG.mem_23_1 ), .C(FIFO_CLK_c), .D(n6335));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2246_2247 (.Q(\REG.mem_23_0 ), .C(FIFO_CLK_c), .D(n6334));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2243_2244 (.Q(\REG.mem_22_31 ), .C(FIFO_CLK_c), .D(n6333));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2240_2241 (.Q(\REG.mem_22_30 ), .C(FIFO_CLK_c), .D(n6332));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2237_2238 (.Q(\REG.mem_22_29 ), .C(FIFO_CLK_c), .D(n6331));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2234_2235 (.Q(\REG.mem_22_28 ), .C(FIFO_CLK_c), .D(n6330));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2231_2232 (.Q(\REG.mem_22_27 ), .C(FIFO_CLK_c), .D(n6329));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2228_2229 (.Q(\REG.mem_22_26 ), .C(FIFO_CLK_c), .D(n6328));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2225_2226 (.Q(\REG.mem_22_25 ), .C(FIFO_CLK_c), .D(n6327));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2222_2223 (.Q(\REG.mem_22_24 ), .C(FIFO_CLK_c), .D(n6326));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2219_2220 (.Q(\REG.mem_22_23 ), .C(FIFO_CLK_c), .D(n6325));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2216_2217 (.Q(\REG.mem_22_22 ), .C(FIFO_CLK_c), .D(n6324));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2213_2214 (.Q(\REG.mem_22_21 ), .C(FIFO_CLK_c), .D(n6323));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2210_2211 (.Q(\REG.mem_22_20 ), .C(FIFO_CLK_c), .D(n6322));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2207_2208 (.Q(\REG.mem_22_19 ), .C(FIFO_CLK_c), .D(n6321));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2204_2205 (.Q(\REG.mem_22_18 ), .C(FIFO_CLK_c), .D(n6320));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2201_2202 (.Q(\REG.mem_22_17 ), .C(FIFO_CLK_c), .D(n6319));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2198_2199 (.Q(\REG.mem_22_16 ), .C(FIFO_CLK_c), .D(n6318));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2195_2196 (.Q(\REG.mem_22_15 ), .C(FIFO_CLK_c), .D(n6317));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2192_2193 (.Q(\REG.mem_22_14 ), .C(FIFO_CLK_c), .D(n6316));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2189_2190 (.Q(\REG.mem_22_13 ), .C(FIFO_CLK_c), .D(n6315));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2186_2187 (.Q(\REG.mem_22_12 ), .C(FIFO_CLK_c), .D(n6314));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2183_2184 (.Q(\REG.mem_22_11 ), .C(FIFO_CLK_c), .D(n6313));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2180_2181 (.Q(\REG.mem_22_10 ), .C(FIFO_CLK_c), .D(n6312));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2177_2178 (.Q(\REG.mem_22_9 ), .C(FIFO_CLK_c), .D(n6311));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2174_2175 (.Q(\REG.mem_22_8 ), .C(FIFO_CLK_c), .D(n6310));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2171_2172 (.Q(\REG.mem_22_7 ), .C(FIFO_CLK_c), .D(n6309));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2168_2169 (.Q(\REG.mem_22_6 ), .C(FIFO_CLK_c), .D(n6308));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2165_2166 (.Q(\REG.mem_22_5 ), .C(FIFO_CLK_c), .D(n6307));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2162_2163 (.Q(\REG.mem_22_4 ), .C(FIFO_CLK_c), .D(n6306));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2159_2160 (.Q(\REG.mem_22_3 ), .C(FIFO_CLK_c), .D(n6305));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2156_2157 (.Q(\REG.mem_22_2 ), .C(FIFO_CLK_c), .D(n6304));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2153_2154 (.Q(\REG.mem_22_1 ), .C(FIFO_CLK_c), .D(n6303));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2150_2151 (.Q(\REG.mem_22_0 ), .C(FIFO_CLK_c), .D(n6302));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2147_2148 (.Q(\REG.mem_21_31 ), .C(FIFO_CLK_c), .D(n6301));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2144_2145 (.Q(\REG.mem_21_30 ), .C(FIFO_CLK_c), .D(n6300));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2141_2142 (.Q(\REG.mem_21_29 ), .C(FIFO_CLK_c), .D(n6299));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2138_2139 (.Q(\REG.mem_21_28 ), .C(FIFO_CLK_c), .D(n6298));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2135_2136 (.Q(\REG.mem_21_27 ), .C(FIFO_CLK_c), .D(n6297));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2132_2133 (.Q(\REG.mem_21_26 ), .C(FIFO_CLK_c), .D(n6296));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2129_2130 (.Q(\REG.mem_21_25 ), .C(FIFO_CLK_c), .D(n6295));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2126_2127 (.Q(\REG.mem_21_24 ), .C(FIFO_CLK_c), .D(n6294));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2123_2124 (.Q(\REG.mem_21_23 ), .C(FIFO_CLK_c), .D(n6293));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2120_2121 (.Q(\REG.mem_21_22 ), .C(FIFO_CLK_c), .D(n6292));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2117_2118 (.Q(\REG.mem_21_21 ), .C(FIFO_CLK_c), .D(n6291));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2114_2115 (.Q(\REG.mem_21_20 ), .C(FIFO_CLK_c), .D(n6290));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2111_2112 (.Q(\REG.mem_21_19 ), .C(FIFO_CLK_c), .D(n6289));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2108_2109 (.Q(\REG.mem_21_18 ), .C(FIFO_CLK_c), .D(n6288));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2105_2106 (.Q(\REG.mem_21_17 ), .C(FIFO_CLK_c), .D(n6287));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2102_2103 (.Q(\REG.mem_21_16 ), .C(FIFO_CLK_c), .D(n6286));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2099_2100 (.Q(\REG.mem_21_15 ), .C(FIFO_CLK_c), .D(n6285));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2096_2097 (.Q(\REG.mem_21_14 ), .C(FIFO_CLK_c), .D(n6284));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2093_2094 (.Q(\REG.mem_21_13 ), .C(FIFO_CLK_c), .D(n6283));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2090_2091 (.Q(\REG.mem_21_12 ), .C(FIFO_CLK_c), .D(n6282));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2087_2088 (.Q(\REG.mem_21_11 ), .C(FIFO_CLK_c), .D(n6281));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2084_2085 (.Q(\REG.mem_21_10 ), .C(FIFO_CLK_c), .D(n6280));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2081_2082 (.Q(\REG.mem_21_9 ), .C(FIFO_CLK_c), .D(n6279));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2078_2079 (.Q(\REG.mem_21_8 ), .C(FIFO_CLK_c), .D(n6278));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2075_2076 (.Q(\REG.mem_21_7 ), .C(FIFO_CLK_c), .D(n6277));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2072_2073 (.Q(\REG.mem_21_6 ), .C(FIFO_CLK_c), .D(n6276));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2069_2070 (.Q(\REG.mem_21_5 ), .C(FIFO_CLK_c), .D(n6275));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2066_2067 (.Q(\REG.mem_21_4 ), .C(FIFO_CLK_c), .D(n6274));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2063_2064 (.Q(\REG.mem_21_3 ), .C(FIFO_CLK_c), .D(n6273));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2060_2061 (.Q(\REG.mem_21_2 ), .C(FIFO_CLK_c), .D(n6272));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2057_2058 (.Q(\REG.mem_21_1 ), .C(FIFO_CLK_c), .D(n6271));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2054_2055 (.Q(\REG.mem_21_0 ), .C(FIFO_CLK_c), .D(n6270));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2051_2052 (.Q(\REG.mem_20_31 ), .C(FIFO_CLK_c), .D(n6269));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2048_2049 (.Q(\REG.mem_20_30 ), .C(FIFO_CLK_c), .D(n6268));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2045_2046 (.Q(\REG.mem_20_29 ), .C(FIFO_CLK_c), .D(n6267));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2042_2043 (.Q(\REG.mem_20_28 ), .C(FIFO_CLK_c), .D(n6266));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2039_2040 (.Q(\REG.mem_20_27 ), .C(FIFO_CLK_c), .D(n6265));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2036_2037 (.Q(\REG.mem_20_26 ), .C(FIFO_CLK_c), .D(n6264));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2033_2034 (.Q(\REG.mem_20_25 ), .C(FIFO_CLK_c), .D(n6263));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2030_2031 (.Q(\REG.mem_20_24 ), .C(FIFO_CLK_c), .D(n6262));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2027_2028 (.Q(\REG.mem_20_23 ), .C(FIFO_CLK_c), .D(n6261));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2024_2025 (.Q(\REG.mem_20_22 ), .C(FIFO_CLK_c), .D(n6260));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2021_2022 (.Q(\REG.mem_20_21 ), .C(FIFO_CLK_c), .D(n6259));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2018_2019 (.Q(\REG.mem_20_20 ), .C(FIFO_CLK_c), .D(n6258));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2015_2016 (.Q(\REG.mem_20_19 ), .C(FIFO_CLK_c), .D(n6257));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2012_2013 (.Q(\REG.mem_20_18 ), .C(FIFO_CLK_c), .D(n6256));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2009_2010 (.Q(\REG.mem_20_17 ), .C(FIFO_CLK_c), .D(n6255));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2006_2007 (.Q(\REG.mem_20_16 ), .C(FIFO_CLK_c), .D(n6254));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2003_2004 (.Q(\REG.mem_20_15 ), .C(FIFO_CLK_c), .D(n6253));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2000_2001 (.Q(\REG.mem_20_14 ), .C(FIFO_CLK_c), .D(n6252));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1997_1998 (.Q(\REG.mem_20_13 ), .C(FIFO_CLK_c), .D(n6251));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1994_1995 (.Q(\REG.mem_20_12 ), .C(FIFO_CLK_c), .D(n6250));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1991_1992 (.Q(\REG.mem_20_11 ), .C(FIFO_CLK_c), .D(n6249));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1988_1989 (.Q(\REG.mem_20_10 ), .C(FIFO_CLK_c), .D(n6248));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1985_1986 (.Q(\REG.mem_20_9 ), .C(FIFO_CLK_c), .D(n6247));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1982_1983 (.Q(\REG.mem_20_8 ), .C(FIFO_CLK_c), .D(n6246));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1979_1980 (.Q(\REG.mem_20_7 ), .C(FIFO_CLK_c), .D(n6245));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1976_1977 (.Q(\REG.mem_20_6 ), .C(FIFO_CLK_c), .D(n6244));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1973_1974 (.Q(\REG.mem_20_5 ), .C(FIFO_CLK_c), .D(n6243));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1970_1971 (.Q(\REG.mem_20_4 ), .C(FIFO_CLK_c), .D(n6242));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1967_1968 (.Q(\REG.mem_20_3 ), .C(FIFO_CLK_c), .D(n6241));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1964_1965 (.Q(\REG.mem_20_2 ), .C(FIFO_CLK_c), .D(n6240));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1961_1962 (.Q(\REG.mem_20_1 ), .C(FIFO_CLK_c), .D(n6239));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1958_1959 (.Q(\REG.mem_20_0 ), .C(FIFO_CLK_c), .D(n6238));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1955_1956 (.Q(\REG.mem_19_31 ), .C(FIFO_CLK_c), .D(n6237));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1952_1953 (.Q(\REG.mem_19_30 ), .C(FIFO_CLK_c), .D(n6236));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1949_1950 (.Q(\REG.mem_19_29 ), .C(FIFO_CLK_c), .D(n6235));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1946_1947 (.Q(\REG.mem_19_28 ), .C(FIFO_CLK_c), .D(n6234));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1943_1944 (.Q(\REG.mem_19_27 ), .C(FIFO_CLK_c), .D(n6233));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1940_1941 (.Q(\REG.mem_19_26 ), .C(FIFO_CLK_c), .D(n6232));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1937_1938 (.Q(\REG.mem_19_25 ), .C(FIFO_CLK_c), .D(n6231));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1934_1935 (.Q(\REG.mem_19_24 ), .C(FIFO_CLK_c), .D(n6230));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1931_1932 (.Q(\REG.mem_19_23 ), .C(FIFO_CLK_c), .D(n6229));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1928_1929 (.Q(\REG.mem_19_22 ), .C(FIFO_CLK_c), .D(n6228));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1925_1926 (.Q(\REG.mem_19_21 ), .C(FIFO_CLK_c), .D(n6227));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1922_1923 (.Q(\REG.mem_19_20 ), .C(FIFO_CLK_c), .D(n6226));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1919_1920 (.Q(\REG.mem_19_19 ), .C(FIFO_CLK_c), .D(n6225));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1916_1917 (.Q(\REG.mem_19_18 ), .C(FIFO_CLK_c), .D(n6224));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1913_1914 (.Q(\REG.mem_19_17 ), .C(FIFO_CLK_c), .D(n6223));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1910_1911 (.Q(\REG.mem_19_16 ), .C(FIFO_CLK_c), .D(n6222));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1907_1908 (.Q(\REG.mem_19_15 ), .C(FIFO_CLK_c), .D(n6221));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1904_1905 (.Q(\REG.mem_19_14 ), .C(FIFO_CLK_c), .D(n6220));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1901_1902 (.Q(\REG.mem_19_13 ), .C(FIFO_CLK_c), .D(n6219));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1898_1899 (.Q(\REG.mem_19_12 ), .C(FIFO_CLK_c), .D(n6218));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1895_1896 (.Q(\REG.mem_19_11 ), .C(FIFO_CLK_c), .D(n6217));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1892_1893 (.Q(\REG.mem_19_10 ), .C(FIFO_CLK_c), .D(n6216));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1889_1890 (.Q(\REG.mem_19_9 ), .C(FIFO_CLK_c), .D(n6215));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1886_1887 (.Q(\REG.mem_19_8 ), .C(FIFO_CLK_c), .D(n6214));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1883_1884 (.Q(\REG.mem_19_7 ), .C(FIFO_CLK_c), .D(n6213));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1880_1881 (.Q(\REG.mem_19_6 ), .C(FIFO_CLK_c), .D(n6212));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1877_1878 (.Q(\REG.mem_19_5 ), .C(FIFO_CLK_c), .D(n6211));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1874_1875 (.Q(\REG.mem_19_4 ), .C(FIFO_CLK_c), .D(n6210));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1871_1872 (.Q(\REG.mem_19_3 ), .C(FIFO_CLK_c), .D(n6209));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1868_1869 (.Q(\REG.mem_19_2 ), .C(FIFO_CLK_c), .D(n6208));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1865_1866 (.Q(\REG.mem_19_1 ), .C(FIFO_CLK_c), .D(n6207));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1862_1863 (.Q(\REG.mem_19_0 ), .C(FIFO_CLK_c), .D(n6206));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1859_1860 (.Q(\REG.mem_18_31 ), .C(FIFO_CLK_c), .D(n6205));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1856_1857 (.Q(\REG.mem_18_30 ), .C(FIFO_CLK_c), .D(n6204));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1853_1854 (.Q(\REG.mem_18_29 ), .C(FIFO_CLK_c), .D(n6203));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1850_1851 (.Q(\REG.mem_18_28 ), .C(FIFO_CLK_c), .D(n6202));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1847_1848 (.Q(\REG.mem_18_27 ), .C(FIFO_CLK_c), .D(n6201));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1844_1845 (.Q(\REG.mem_18_26 ), .C(FIFO_CLK_c), .D(n6200));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1841_1842 (.Q(\REG.mem_18_25 ), .C(FIFO_CLK_c), .D(n6199));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1838_1839 (.Q(\REG.mem_18_24 ), .C(FIFO_CLK_c), .D(n6198));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1835_1836 (.Q(\REG.mem_18_23 ), .C(FIFO_CLK_c), .D(n6197));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1832_1833 (.Q(\REG.mem_18_22 ), .C(FIFO_CLK_c), .D(n6196));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1829_1830 (.Q(\REG.mem_18_21 ), .C(FIFO_CLK_c), .D(n6195));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1826_1827 (.Q(\REG.mem_18_20 ), .C(FIFO_CLK_c), .D(n6194));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1823_1824 (.Q(\REG.mem_18_19 ), .C(FIFO_CLK_c), .D(n6193));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1820_1821 (.Q(\REG.mem_18_18 ), .C(FIFO_CLK_c), .D(n6192));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1817_1818 (.Q(\REG.mem_18_17 ), .C(FIFO_CLK_c), .D(n6191));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1814_1815 (.Q(\REG.mem_18_16 ), .C(FIFO_CLK_c), .D(n6190));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1811_1812 (.Q(\REG.mem_18_15 ), .C(FIFO_CLK_c), .D(n6189));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1808_1809 (.Q(\REG.mem_18_14 ), .C(FIFO_CLK_c), .D(n6188));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1805_1806 (.Q(\REG.mem_18_13 ), .C(FIFO_CLK_c), .D(n6187));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1802_1803 (.Q(\REG.mem_18_12 ), .C(FIFO_CLK_c), .D(n6186));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1799_1800 (.Q(\REG.mem_18_11 ), .C(FIFO_CLK_c), .D(n6185));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1796_1797 (.Q(\REG.mem_18_10 ), .C(FIFO_CLK_c), .D(n6184));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1793_1794 (.Q(\REG.mem_18_9 ), .C(FIFO_CLK_c), .D(n6183));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1790_1791 (.Q(\REG.mem_18_8 ), .C(FIFO_CLK_c), .D(n6182));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1787_1788 (.Q(\REG.mem_18_7 ), .C(FIFO_CLK_c), .D(n6181));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1784_1785 (.Q(\REG.mem_18_6 ), .C(FIFO_CLK_c), .D(n6180));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1781_1782 (.Q(\REG.mem_18_5 ), .C(FIFO_CLK_c), .D(n6179));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1778_1779 (.Q(\REG.mem_18_4 ), .C(FIFO_CLK_c), .D(n6178));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1775_1776 (.Q(\REG.mem_18_3 ), .C(FIFO_CLK_c), .D(n6177));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1772_1773 (.Q(\REG.mem_18_2 ), .C(FIFO_CLK_c), .D(n6176));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1769_1770 (.Q(\REG.mem_18_1 ), .C(FIFO_CLK_c), .D(n6175));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1766_1767 (.Q(\REG.mem_18_0 ), .C(FIFO_CLK_c), .D(n6174));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1763_1764 (.Q(\REG.mem_17_31 ), .C(FIFO_CLK_c), .D(n6173));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1760_1761 (.Q(\REG.mem_17_30 ), .C(FIFO_CLK_c), .D(n6172));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1757_1758 (.Q(\REG.mem_17_29 ), .C(FIFO_CLK_c), .D(n6171));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1754_1755 (.Q(\REG.mem_17_28 ), .C(FIFO_CLK_c), .D(n6170));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1751_1752 (.Q(\REG.mem_17_27 ), .C(FIFO_CLK_c), .D(n6169));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1748_1749 (.Q(\REG.mem_17_26 ), .C(FIFO_CLK_c), .D(n6168));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1745_1746 (.Q(\REG.mem_17_25 ), .C(FIFO_CLK_c), .D(n6167));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1742_1743 (.Q(\REG.mem_17_24 ), .C(FIFO_CLK_c), .D(n6166));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1739_1740 (.Q(\REG.mem_17_23 ), .C(FIFO_CLK_c), .D(n6165));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1736_1737 (.Q(\REG.mem_17_22 ), .C(FIFO_CLK_c), .D(n6164));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1733_1734 (.Q(\REG.mem_17_21 ), .C(FIFO_CLK_c), .D(n6163));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1730_1731 (.Q(\REG.mem_17_20 ), .C(FIFO_CLK_c), .D(n6162));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1727_1728 (.Q(\REG.mem_17_19 ), .C(FIFO_CLK_c), .D(n6161));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1724_1725 (.Q(\REG.mem_17_18 ), .C(FIFO_CLK_c), .D(n6160));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1721_1722 (.Q(\REG.mem_17_17 ), .C(FIFO_CLK_c), .D(n6159));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1718_1719 (.Q(\REG.mem_17_16 ), .C(FIFO_CLK_c), .D(n6158));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1715_1716 (.Q(\REG.mem_17_15 ), .C(FIFO_CLK_c), .D(n6157));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1712_1713 (.Q(\REG.mem_17_14 ), .C(FIFO_CLK_c), .D(n6156));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1709_1710 (.Q(\REG.mem_17_13 ), .C(FIFO_CLK_c), .D(n6155));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1706_1707 (.Q(\REG.mem_17_12 ), .C(FIFO_CLK_c), .D(n6154));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1703_1704 (.Q(\REG.mem_17_11 ), .C(FIFO_CLK_c), .D(n6153));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1700_1701 (.Q(\REG.mem_17_10 ), .C(FIFO_CLK_c), .D(n6152));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1697_1698 (.Q(\REG.mem_17_9 ), .C(FIFO_CLK_c), .D(n6151));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1694_1695 (.Q(\REG.mem_17_8 ), .C(FIFO_CLK_c), .D(n6150));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1691_1692 (.Q(\REG.mem_17_7 ), .C(FIFO_CLK_c), .D(n6149));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1688_1689 (.Q(\REG.mem_17_6 ), .C(FIFO_CLK_c), .D(n6148));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1685_1686 (.Q(\REG.mem_17_5 ), .C(FIFO_CLK_c), .D(n6147));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1682_1683 (.Q(\REG.mem_17_4 ), .C(FIFO_CLK_c), .D(n6146));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1679_1680 (.Q(\REG.mem_17_3 ), .C(FIFO_CLK_c), .D(n6145));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1676_1677 (.Q(\REG.mem_17_2 ), .C(FIFO_CLK_c), .D(n6144));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1673_1674 (.Q(\REG.mem_17_1 ), .C(FIFO_CLK_c), .D(n6143));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1670_1671 (.Q(\REG.mem_17_0 ), .C(FIFO_CLK_c), .D(n6142));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1667_1668 (.Q(\REG.mem_16_31 ), .C(FIFO_CLK_c), .D(n6141));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1664_1665 (.Q(\REG.mem_16_30 ), .C(FIFO_CLK_c), .D(n6140));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1661_1662 (.Q(\REG.mem_16_29 ), .C(FIFO_CLK_c), .D(n6139));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1658_1659 (.Q(\REG.mem_16_28 ), .C(FIFO_CLK_c), .D(n6138));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1655_1656 (.Q(\REG.mem_16_27 ), .C(FIFO_CLK_c), .D(n6137));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1652_1653 (.Q(\REG.mem_16_26 ), .C(FIFO_CLK_c), .D(n6136));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1649_1650 (.Q(\REG.mem_16_25 ), .C(FIFO_CLK_c), .D(n6135));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1646_1647 (.Q(\REG.mem_16_24 ), .C(FIFO_CLK_c), .D(n6134));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1643_1644 (.Q(\REG.mem_16_23 ), .C(FIFO_CLK_c), .D(n6133));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1640_1641 (.Q(\REG.mem_16_22 ), .C(FIFO_CLK_c), .D(n6132));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1637_1638 (.Q(\REG.mem_16_21 ), .C(FIFO_CLK_c), .D(n6131));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1634_1635 (.Q(\REG.mem_16_20 ), .C(FIFO_CLK_c), .D(n6130));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1631_1632 (.Q(\REG.mem_16_19 ), .C(FIFO_CLK_c), .D(n6129));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1628_1629 (.Q(\REG.mem_16_18 ), .C(FIFO_CLK_c), .D(n6128));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1625_1626 (.Q(\REG.mem_16_17 ), .C(FIFO_CLK_c), .D(n6127));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1622_1623 (.Q(\REG.mem_16_16 ), .C(FIFO_CLK_c), .D(n6126));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1619_1620 (.Q(\REG.mem_16_15 ), .C(FIFO_CLK_c), .D(n6125));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1616_1617 (.Q(\REG.mem_16_14 ), .C(FIFO_CLK_c), .D(n6124));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1613_1614 (.Q(\REG.mem_16_13 ), .C(FIFO_CLK_c), .D(n6123));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1610_1611 (.Q(\REG.mem_16_12 ), .C(FIFO_CLK_c), .D(n6122));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1607_1608 (.Q(\REG.mem_16_11 ), .C(FIFO_CLK_c), .D(n6121));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1604_1605 (.Q(\REG.mem_16_10 ), .C(FIFO_CLK_c), .D(n6120));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1601_1602 (.Q(\REG.mem_16_9 ), .C(FIFO_CLK_c), .D(n6119));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1598_1599 (.Q(\REG.mem_16_8 ), .C(FIFO_CLK_c), .D(n6118));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1595_1596 (.Q(\REG.mem_16_7 ), .C(FIFO_CLK_c), .D(n6117));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1592_1593 (.Q(\REG.mem_16_6 ), .C(FIFO_CLK_c), .D(n6116));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1589_1590 (.Q(\REG.mem_16_5 ), .C(FIFO_CLK_c), .D(n6115));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1586_1587 (.Q(\REG.mem_16_4 ), .C(FIFO_CLK_c), .D(n6114));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1583_1584 (.Q(\REG.mem_16_3 ), .C(FIFO_CLK_c), .D(n6113));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1580_1581 (.Q(\REG.mem_16_2 ), .C(FIFO_CLK_c), .D(n6112));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1577_1578 (.Q(\REG.mem_16_1 ), .C(FIFO_CLK_c), .D(n6111));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1574_1575 (.Q(\REG.mem_16_0 ), .C(FIFO_CLK_c), .D(n6110));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1571_1572 (.Q(\REG.mem_15_31 ), .C(FIFO_CLK_c), .D(n6109));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1568_1569 (.Q(\REG.mem_15_30 ), .C(FIFO_CLK_c), .D(n6108));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1565_1566 (.Q(\REG.mem_15_29 ), .C(FIFO_CLK_c), .D(n6107));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1562_1563 (.Q(\REG.mem_15_28 ), .C(FIFO_CLK_c), .D(n6106));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1559_1560 (.Q(\REG.mem_15_27 ), .C(FIFO_CLK_c), .D(n6105));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1556_1557 (.Q(\REG.mem_15_26 ), .C(FIFO_CLK_c), .D(n6104));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1553_1554 (.Q(\REG.mem_15_25 ), .C(FIFO_CLK_c), .D(n6103));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1550_1551 (.Q(\REG.mem_15_24 ), .C(FIFO_CLK_c), .D(n6102));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1547_1548 (.Q(\REG.mem_15_23 ), .C(FIFO_CLK_c), .D(n6101));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1544_1545 (.Q(\REG.mem_15_22 ), .C(FIFO_CLK_c), .D(n6100));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1541_1542 (.Q(\REG.mem_15_21 ), .C(FIFO_CLK_c), .D(n6099));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1538_1539 (.Q(\REG.mem_15_20 ), .C(FIFO_CLK_c), .D(n6098));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1535_1536 (.Q(\REG.mem_15_19 ), .C(FIFO_CLK_c), .D(n6097));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1532_1533 (.Q(\REG.mem_15_18 ), .C(FIFO_CLK_c), .D(n6096));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1529_1530 (.Q(\REG.mem_15_17 ), .C(FIFO_CLK_c), .D(n6095));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1526_1527 (.Q(\REG.mem_15_16 ), .C(FIFO_CLK_c), .D(n6094));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1523_1524 (.Q(\REG.mem_15_15 ), .C(FIFO_CLK_c), .D(n6093));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1520_1521 (.Q(\REG.mem_15_14 ), .C(FIFO_CLK_c), .D(n6092));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1517_1518 (.Q(\REG.mem_15_13 ), .C(FIFO_CLK_c), .D(n6091));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1514_1515 (.Q(\REG.mem_15_12 ), .C(FIFO_CLK_c), .D(n6090));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1511_1512 (.Q(\REG.mem_15_11 ), .C(FIFO_CLK_c), .D(n6089));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1508_1509 (.Q(\REG.mem_15_10 ), .C(FIFO_CLK_c), .D(n6088));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4602_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_14_30 ), .O(n6076));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4602_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1505_1506 (.Q(\REG.mem_15_9 ), .C(FIFO_CLK_c), .D(n6087));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1502_1503 (.Q(\REG.mem_15_8 ), .C(FIFO_CLK_c), .D(n6086));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1499_1500 (.Q(\REG.mem_15_7 ), .C(FIFO_CLK_c), .D(n6085));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1496_1497 (.Q(\REG.mem_15_6 ), .C(FIFO_CLK_c), .D(n6084));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1493_1494 (.Q(\REG.mem_15_5 ), .C(FIFO_CLK_c), .D(n6083));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1490_1491 (.Q(\REG.mem_15_4 ), .C(FIFO_CLK_c), .D(n6082));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1487_1488 (.Q(\REG.mem_15_3 ), .C(FIFO_CLK_c), .D(n6081));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1484_1485 (.Q(\REG.mem_15_2 ), .C(FIFO_CLK_c), .D(n6080));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1481_1482 (.Q(\REG.mem_15_1 ), .C(FIFO_CLK_c), .D(n6079));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1478_1479 (.Q(\REG.mem_15_0 ), .C(FIFO_CLK_c), .D(n6078));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12772 (.I0(rd_addr_r[1]), .I1(n13354), 
            .I2(n13355), .I3(rd_addr_r[2]), .O(n14953));
    defparam rd_addr_r_1__bdd_4_lut_12772.LUT_INIT = 16'he4aa;
    SB_DFF i1475_1476 (.Q(\REG.mem_14_31 ), .C(FIFO_CLK_c), .D(n6077));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1472_1473 (.Q(\REG.mem_14_30 ), .C(FIFO_CLK_c), .D(n6076));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1469_1470 (.Q(\REG.mem_14_29 ), .C(FIFO_CLK_c), .D(n6075));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1466_1467 (.Q(\REG.mem_14_28 ), .C(FIFO_CLK_c), .D(n6074));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1463_1464 (.Q(\REG.mem_14_27 ), .C(FIFO_CLK_c), .D(n6073));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1460_1461 (.Q(\REG.mem_14_26 ), .C(FIFO_CLK_c), .D(n6072));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1457_1458 (.Q(\REG.mem_14_25 ), .C(FIFO_CLK_c), .D(n6071));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1454_1455 (.Q(\REG.mem_14_24 ), .C(FIFO_CLK_c), .D(n6070));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i320_321 (.Q(\REG.mem_2_30 ), .C(FIFO_CLK_c), .D(n5692));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14953_bdd_4_lut (.I0(n14953), .I1(n13352), .I2(n13351), .I3(rd_addr_r[2]), 
            .O(n14956));
    defparam n14953_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15637_bdd_4_lut (.I0(n15637), .I1(\REG.mem_5_30 ), .I2(\REG.mem_4_30 ), 
            .I3(rd_addr_r[1]), .O(n15640));
    defparam n15637_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12767 (.I0(rd_addr_r[3]), .I1(n13483), 
            .I2(n13484), .I3(rd_addr_r[4]), .O(n14947));
    defparam rd_addr_r_3__bdd_4_lut_12767.LUT_INIT = 16'he4aa;
    SB_LUT4 n14947_bdd_4_lut (.I0(n14947), .I1(n13379), .I2(n14938), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[2]));
    defparam n14947_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i317_318 (.Q(\REG.mem_2_29 ), .C(FIFO_CLK_c), .D(n5691));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_13396 (.I0(rd_addr_r[3]), .I1(n13741), 
            .I2(n13742), .I3(rd_addr_r[4]), .O(n15631));
    defparam rd_addr_r_3__bdd_4_lut_13396.LUT_INIT = 16'he4aa;
    SB_DFF i314_315 (.Q(\REG.mem_2_28 ), .C(FIFO_CLK_c), .D(n5690));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n15631_bdd_4_lut (.I0(n15631), .I1(n13685), .I2(n15472), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[15]));
    defparam n15631_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4601_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_14_29 ), .O(n6075));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4601_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12762 (.I0(rd_addr_r[1]), .I1(n13144), 
            .I2(n13145), .I3(rd_addr_r[2]), .O(n14941));
    defparam rd_addr_r_1__bdd_4_lut_12762.LUT_INIT = 16'he4aa;
    SB_LUT4 n14941_bdd_4_lut (.I0(n14941), .I1(n13088), .I2(n13087), .I3(rd_addr_r[2]), 
            .O(n14944));
    defparam n14941_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12752 (.I0(rd_addr_r[1]), .I1(n13342), 
            .I2(n13343), .I3(rd_addr_r[2]), .O(n14935));
    defparam rd_addr_r_1__bdd_4_lut_12752.LUT_INIT = 16'he4aa;
    SB_DFF i1451_1452 (.Q(\REG.mem_14_23 ), .C(FIFO_CLK_c), .D(n6069));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i11271_3_lut (.I0(n14548), .I1(n15808), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13382));
    defparam i11271_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1448_1449 (.Q(\REG.mem_14_22 ), .C(FIFO_CLK_c), .D(n6068));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1445_1446 (.Q(\REG.mem_14_21 ), .C(FIFO_CLK_c), .D(n6067));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1442_1443 (.Q(\REG.mem_14_20 ), .C(FIFO_CLK_c), .D(n6066));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1439_1440 (.Q(\REG.mem_14_19 ), .C(FIFO_CLK_c), .D(n6065));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1436_1437 (.Q(\REG.mem_14_18 ), .C(FIFO_CLK_c), .D(n6064));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1433_1434 (.Q(\REG.mem_14_17 ), .C(FIFO_CLK_c), .D(n6063));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1430_1431 (.Q(\REG.mem_14_16 ), .C(FIFO_CLK_c), .D(n6062));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1427_1428 (.Q(\REG.mem_14_15 ), .C(FIFO_CLK_c), .D(n6061));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i311_312 (.Q(\REG.mem_2_27 ), .C(FIFO_CLK_c), .D(n5689));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i11273_3_lut (.I0(\REG.mem_0_1 ), .I1(\REG.mem_1_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13384));
    defparam i11273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11274_3_lut (.I0(\REG.mem_2_1 ), .I1(\REG.mem_3_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13385));
    defparam i11274_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n14935_bdd_4_lut (.I0(n14935), .I1(n13340), .I2(n13339), .I3(rd_addr_r[2]), 
            .O(n14938));
    defparam n14935_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i308_309 (.Q(\REG.mem_2_26 ), .C(FIFO_CLK_c), .D(n5688));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12757 (.I0(rd_addr_r[3]), .I1(n14800), 
            .I2(n13157), .I3(rd_addr_r[4]), .O(n14929));
    defparam rd_addr_r_3__bdd_4_lut_12757.LUT_INIT = 16'he4aa;
    SB_DFF i305_306 (.Q(\REG.mem_2_25 ), .C(FIFO_CLK_c), .D(n5687));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1424_1425 (.Q(\REG.mem_14_14 ), .C(FIFO_CLK_c), .D(n6060));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13371 (.I0(rd_addr_r[1]), .I1(n13795), 
            .I2(n13796), .I3(rd_addr_r[2]), .O(n15625));
    defparam rd_addr_r_1__bdd_4_lut_13371.LUT_INIT = 16'he4aa;
    SB_LUT4 n15625_bdd_4_lut (.I0(n15625), .I1(n13787), .I2(n13786), .I3(rd_addr_r[2]), 
            .O(n15628));
    defparam n15625_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11369_3_lut (.I0(\REG.mem_16_0 ), .I1(\REG.mem_17_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13480));
    defparam i11369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n14929_bdd_4_lut (.I0(n14929), .I1(n13139), .I2(n14746), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[3]));
    defparam n14929_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i30_2_lut (.I0(n14), .I1(wr_addr_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n30));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12483 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_12 ), 
            .I2(\REG.mem_19_12 ), .I3(rd_addr_r[1]), .O(n14611));
    defparam rd_addr_r_0__bdd_4_lut_12483.LUT_INIT = 16'he4aa;
    SB_DFF i1421_1422 (.Q(\REG.mem_14_13 ), .C(FIFO_CLK_c), .D(n6059));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1418_1419 (.Q(\REG.mem_14_12 ), .C(FIFO_CLK_c), .D(n6058));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1415_1416 (.Q(\REG.mem_14_11 ), .C(FIFO_CLK_c), .D(n6057));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1412_1413 (.Q(\REG.mem_14_10 ), .C(FIFO_CLK_c), .D(n6056));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1409_1410 (.Q(\REG.mem_14_9 ), .C(FIFO_CLK_c), .D(n6055));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1406_1407 (.Q(\REG.mem_14_8 ), .C(FIFO_CLK_c), .D(n6054));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1403_1404 (.Q(\REG.mem_14_7 ), .C(FIFO_CLK_c), .D(n6053));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14611_bdd_4_lut (.I0(n14611), .I1(\REG.mem_17_12 ), .I2(\REG.mem_16_12 ), 
            .I3(rd_addr_r[1]), .O(n14614));
    defparam n14611_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i302_303 (.Q(\REG.mem_2_24 ), .C(FIFO_CLK_c), .D(n5686));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i11370_3_lut (.I0(\REG.mem_18_0 ), .I1(\REG.mem_19_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13481));
    defparam i11370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11277_3_lut (.I0(\REG.mem_6_1 ), .I1(\REG.mem_7_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13388));
    defparam i11277_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i299_300 (.Q(\REG.mem_2_23 ), .C(FIFO_CLK_c), .D(n5685));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i11276_3_lut (.I0(\REG.mem_4_1 ), .I1(\REG.mem_5_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13387));
    defparam i11276_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1400_1401 (.Q(\REG.mem_14_6 ), .C(FIFO_CLK_c), .D(n6052));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1397_1398 (.Q(\REG.mem_14_5 ), .C(FIFO_CLK_c), .D(n6051));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1394_1395 (.Q(\REG.mem_14_4 ), .C(FIFO_CLK_c), .D(n6050));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1391_1392 (.Q(\REG.mem_14_3 ), .C(FIFO_CLK_c), .D(n6049));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1388_1389 (.Q(\REG.mem_14_2 ), .C(FIFO_CLK_c), .D(n6048));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1385_1386 (.Q(\REG.mem_14_1 ), .C(FIFO_CLK_c), .D(n6047));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1382_1383 (.Q(\REG.mem_14_0 ), .C(FIFO_CLK_c), .D(n6046));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1379_1380 (.Q(\REG.mem_13_31 ), .C(FIFO_CLK_c), .D(n6045));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i11382_3_lut (.I0(\REG.mem_22_0 ), .I1(\REG.mem_23_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13493));
    defparam i11382_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1376_1377 (.Q(\REG.mem_13_30 ), .C(FIFO_CLK_c), .D(n6044));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i11381_3_lut (.I0(\REG.mem_20_0 ), .I1(\REG.mem_21_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13492));
    defparam i11381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13331 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_21 ), 
            .I2(\REG.mem_7_21 ), .I3(rd_addr_r[1]), .O(n15613));
    defparam rd_addr_r_0__bdd_4_lut_13331.LUT_INIT = 16'he4aa;
    SB_LUT4 n15613_bdd_4_lut (.I0(n15613), .I1(\REG.mem_5_21 ), .I2(\REG.mem_4_21 ), 
            .I3(rd_addr_r[1]), .O(n15616));
    defparam n15613_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4600_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_14_28 ), .O(n6074));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4600_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12827 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_5 ), 
            .I2(\REG.mem_19_5 ), .I3(rd_addr_r[1]), .O(n14923));
    defparam rd_addr_r_0__bdd_4_lut_12827.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_13656 (.I0(rd_addr_r[2]), .I1(n13764), 
            .I2(n13668), .I3(rd_addr_r[3]), .O(n15607));
    defparam rd_addr_r_2__bdd_4_lut_13656.LUT_INIT = 16'he4aa;
    SB_LUT4 i4599_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_14_27 ), .O(n6073));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4599_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1373_1374 (.Q(\REG.mem_13_29 ), .C(FIFO_CLK_c), .D(n6043));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n15607_bdd_4_lut (.I0(n15607), .I1(n13761), .I2(n13683), .I3(rd_addr_r[3]), 
            .O(n15610));
    defparam n15607_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4598_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_14_26 ), .O(n6072));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4598_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4597_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_14_25 ), .O(n6071));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4597_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1370_1371 (.Q(\REG.mem_13_28 ), .C(FIFO_CLK_c), .D(n6042));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14923_bdd_4_lut (.I0(n14923), .I1(\REG.mem_17_5 ), .I2(\REG.mem_16_5 ), 
            .I3(rd_addr_r[1]), .O(n14926));
    defparam n14923_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4596_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_14_24 ), .O(n6070));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4596_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4595_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_14_23 ), .O(n6069));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4595_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1367_1368 (.Q(\REG.mem_13_27 ), .C(FIFO_CLK_c), .D(n6041));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1364_1365 (.Q(\REG.mem_13_26 ), .C(FIFO_CLK_c), .D(n6040));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1361_1362 (.Q(\REG.mem_13_25 ), .C(FIFO_CLK_c), .D(n6039));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1358_1359 (.Q(\REG.mem_13_24 ), .C(FIFO_CLK_c), .D(n6038));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4594_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_14_22 ), .O(n6068));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4594_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1355_1356 (.Q(\REG.mem_13_23 ), .C(FIFO_CLK_c), .D(n6037));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1352_1353 (.Q(\REG.mem_13_22 ), .C(FIFO_CLK_c), .D(n6036));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1349_1350 (.Q(\REG.mem_13_21 ), .C(FIFO_CLK_c), .D(n6035));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1346_1347 (.Q(\REG.mem_13_20 ), .C(FIFO_CLK_c), .D(n6034));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1343_1344 (.Q(\REG.mem_13_19 ), .C(FIFO_CLK_c), .D(n6033));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1340_1341 (.Q(\REG.mem_13_18 ), .C(FIFO_CLK_c), .D(n6032));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4593_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_14_21 ), .O(n6067));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4593_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1337_1338 (.Q(\REG.mem_13_17 ), .C(FIFO_CLK_c), .D(n6031));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1334_1335 (.Q(\REG.mem_13_16 ), .C(FIFO_CLK_c), .D(n6030));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1331_1332 (.Q(\REG.mem_13_15 ), .C(FIFO_CLK_c), .D(n6029));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1328_1329 (.Q(\REG.mem_13_14 ), .C(FIFO_CLK_c), .D(n6028));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4592_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_14_20 ), .O(n6066));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4592_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4591_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_14_19 ), .O(n6065));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4591_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1325_1326 (.Q(\REG.mem_13_13 ), .C(FIFO_CLK_c), .D(n6027));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1322_1323 (.Q(\REG.mem_13_12 ), .C(FIFO_CLK_c), .D(n6026));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12777 (.I0(rd_addr_r[2]), .I1(n13989), 
            .I2(n13614), .I3(rd_addr_r[3]), .O(n14917));
    defparam rd_addr_r_2__bdd_4_lut_12777.LUT_INIT = 16'he4aa;
    SB_DFF i1319_1320 (.Q(\REG.mem_13_11 ), .C(FIFO_CLK_c), .D(n6025));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1316_1317 (.Q(\REG.mem_13_10 ), .C(FIFO_CLK_c), .D(n6024));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1313_1314 (.Q(\REG.mem_13_9 ), .C(FIFO_CLK_c), .D(n6023));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1310_1311 (.Q(\REG.mem_13_8 ), .C(FIFO_CLK_c), .D(n6022));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1307_1308 (.Q(\REG.mem_13_7 ), .C(FIFO_CLK_c), .D(n6021));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i296_297 (.Q(\REG.mem_2_22 ), .C(FIFO_CLK_c), .D(n5684));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1304_1305 (.Q(\REG.mem_13_6 ), .C(FIFO_CLK_c), .D(n6020));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1301_1302 (.Q(\REG.mem_13_5 ), .C(FIFO_CLK_c), .D(n6019));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1298_1299 (.Q(\REG.mem_13_4 ), .C(FIFO_CLK_c), .D(n6018));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13311 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_28 ), 
            .I2(\REG.mem_15_28 ), .I3(rd_addr_r[1]), .O(n15601));
    defparam rd_addr_r_0__bdd_4_lut_13311.LUT_INIT = 16'he4aa;
    SB_LUT4 n15601_bdd_4_lut (.I0(n15601), .I1(\REG.mem_13_28 ), .I2(\REG.mem_12_28 ), 
            .I3(rd_addr_r[1]), .O(n15604));
    defparam n15601_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14917_bdd_4_lut (.I0(n14917), .I1(n13983), .I2(n13629), .I3(rd_addr_r[3]), 
            .O(n14920));
    defparam n14917_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1295_1296 (.Q(\REG.mem_13_3 ), .C(FIFO_CLK_c), .D(n6017));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12737 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_5 ), 
            .I2(\REG.mem_23_5 ), .I3(rd_addr_r[1]), .O(n14911));
    defparam rd_addr_r_0__bdd_4_lut_12737.LUT_INIT = 16'he4aa;
    SB_DFF i1292_1293 (.Q(\REG.mem_13_2 ), .C(FIFO_CLK_c), .D(n6016));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4590_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_14_18 ), .O(n6064));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4590_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4589_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_14_17 ), .O(n6063));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4589_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i293_294 (.Q(\REG.mem_2_21 ), .C(FIFO_CLK_c), .D(n5683));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1289_1290 (.Q(\REG.mem_13_1 ), .C(FIFO_CLK_c), .D(n6015));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i290_291 (.Q(\REG.mem_2_20 ), .C(FIFO_CLK_c), .D(n5682));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14911_bdd_4_lut (.I0(n14911), .I1(\REG.mem_21_5 ), .I2(\REG.mem_20_5 ), 
            .I3(rd_addr_r[1]), .O(n14914));
    defparam n14911_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13301 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_10 ), 
            .I2(\REG.mem_31_10 ), .I3(rd_addr_r[1]), .O(n15595));
    defparam rd_addr_r_0__bdd_4_lut_13301.LUT_INIT = 16'he4aa;
    SB_DFF i1286_1287 (.Q(\REG.mem_13_0 ), .C(FIFO_CLK_c), .D(n6014));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n15595_bdd_4_lut (.I0(n15595), .I1(\REG.mem_29_10 ), .I2(\REG.mem_28_10 ), 
            .I3(rd_addr_r[1]), .O(n15598));
    defparam n15595_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i287_288 (.Q(\REG.mem_2_19 ), .C(FIFO_CLK_c), .D(n5681));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1283_1284 (.Q(\REG.mem_12_31 ), .C(FIFO_CLK_c), .D(n6013));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4588_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_14_16 ), .O(n6062));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4588_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rp_sync2_r_5__I_0_124_i1_2_lut (.I0(rp_sync2_r[4]), .I1(rp_sync2_r[5]), 
            .I2(GND_net), .I3(GND_net), .O(rp_sync_w[4]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam rp_sync2_r_5__I_0_124_i1_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i4587_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_14_15 ), .O(n6061));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4587_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut (.I0(rp_sync2_r[2]), .I1(rp_sync_w[3]), .I2(GND_net), 
            .I3(GND_net), .O(rp_sync_w[2]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFF i1280_1281 (.Q(\REG.mem_12_30 ), .C(FIFO_CLK_c), .D(n6012));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1277_1278 (.Q(\REG.mem_12_29 ), .C(FIFO_CLK_c), .D(n6011));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4586_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_14_14 ), .O(n6060));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4586_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4585_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_14_13 ), .O(n6059));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4585_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4584_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_14_12 ), .O(n6058));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4584_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12727 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_30 ), 
            .I2(\REG.mem_3_30 ), .I3(rd_addr_r[1]), .O(n14899));
    defparam rd_addr_r_0__bdd_4_lut_12727.LUT_INIT = 16'he4aa;
    SB_LUT4 i4583_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_14_11 ), .O(n6057));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4583_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1274_1275 (.Q(\REG.mem_12_28 ), .C(FIFO_CLK_c), .D(n6010));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4582_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_14_10 ), .O(n6056));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4582_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14899_bdd_4_lut (.I0(n14899), .I1(\REG.mem_1_30 ), .I2(\REG.mem_0_30 ), 
            .I3(rd_addr_r[1]), .O(n14902));
    defparam n14899_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4581_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_14_9 ), .O(n6055));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4581_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i284_285 (.Q(\REG.mem_2_18 ), .C(FIFO_CLK_c), .D(n5680));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12717 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_19 ), 
            .I2(\REG.mem_3_19 ), .I3(rd_addr_r[1]), .O(n14893));
    defparam rd_addr_r_0__bdd_4_lut_12717.LUT_INIT = 16'he4aa;
    SB_LUT4 i4580_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_14_8 ), .O(n6054));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4580_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13296 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_21 ), 
            .I2(\REG.mem_11_21 ), .I3(rd_addr_r[1]), .O(n15583));
    defparam rd_addr_r_0__bdd_4_lut_13296.LUT_INIT = 16'he4aa;
    SB_LUT4 i4579_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_14_7 ), .O(n6053));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4579_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4578_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_14_6 ), .O(n6052));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4578_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12478 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_21 ), 
            .I2(\REG.mem_31_21 ), .I3(rd_addr_r[1]), .O(n14599));
    defparam rd_addr_r_0__bdd_4_lut_12478.LUT_INIT = 16'he4aa;
    SB_LUT4 n14893_bdd_4_lut (.I0(n14893), .I1(\REG.mem_1_19 ), .I2(\REG.mem_0_19 ), 
            .I3(rd_addr_r[1]), .O(n13161));
    defparam n14893_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4088_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_0_4 ), .O(n5562));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4088_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4577_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_14_5 ), .O(n6051));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4577_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i281_282 (.Q(\REG.mem_2_17 ), .C(FIFO_CLK_c), .D(n5679));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1271_1272 (.Q(\REG.mem_12_27 ), .C(FIFO_CLK_c), .D(n6009));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1268_1269 (.Q(\REG.mem_12_26 ), .C(FIFO_CLK_c), .D(n6008));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4576_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_14_4 ), .O(n6050));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4576_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12712 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_19 ), 
            .I2(\REG.mem_7_19 ), .I3(rd_addr_r[1]), .O(n14887));
    defparam rd_addr_r_0__bdd_4_lut_12712.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_68 (.I0(rp_sync2_r[0]), .I1(rp_sync_w[1]), .I2(GND_net), 
            .I3(GND_net), .O(rp_sync_w[0]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_adj_68.LUT_INIT = 16'h6666;
    SB_LUT4 n14887_bdd_4_lut (.I0(n14887), .I1(\REG.mem_5_19 ), .I2(\REG.mem_4_19 ), 
            .I3(rd_addr_r[1]), .O(n13164));
    defparam n14887_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15583_bdd_4_lut (.I0(n15583), .I1(\REG.mem_9_21 ), .I2(\REG.mem_8_21 ), 
            .I3(rd_addr_r[1]), .O(n15586));
    defparam n15583_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut (.I0(rp_sync2_r[3]), .I1(rp_sync2_r[4]), .I2(rp_sync2_r[5]), 
            .I3(GND_net), .O(rp_sync_w[3]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i2_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i4575_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_14_3 ), .O(n6049));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4575_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_4_lut (.I0(wr_addr_p1_w[2]), .I1(wr_addr_p1_w[5]), .I2(rp_sync_w[2]), 
            .I3(rp_sync2_r[5]), .O(n8_adj_1377));
    defparam i2_4_lut.LUT_INIT = 16'h1248;
    SB_DFF i278_279 (.Q(\REG.mem_2_16 ), .C(FIFO_CLK_c), .D(n5678));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10885_4_lut (.I0(wr_addr_p1_w[3]), .I1(\wr_addr_p1_w[0] ), 
            .I2(rp_sync_w[3]), .I3(rp_sync_w[0]), .O(n12994));
    defparam i10885_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 n14599_bdd_4_lut (.I0(n14599), .I1(\REG.mem_29_21 ), .I2(\REG.mem_28_21 ), 
            .I3(rd_addr_r[1]), .O(n14602));
    defparam n14599_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10863_4_lut (.I0(wr_addr_p1_w[4]), .I1(wr_addr_p1_w[1]), .I2(rp_sync_w[4]), 
            .I3(rp_sync_w[1]), .O(n12970));
    defparam i10863_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13286 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_13 ), 
            .I2(\REG.mem_7_13 ), .I3(rd_addr_r[1]), .O(n15571));
    defparam rd_addr_r_0__bdd_4_lut_13286.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12742 (.I0(rd_addr_r[3]), .I1(n14794), 
            .I2(n13154), .I3(rd_addr_r[4]), .O(n14881));
    defparam rd_addr_r_3__bdd_4_lut_12742.LUT_INIT = 16'he4aa;
    SB_DFF i275_276 (.Q(\REG.mem_2_15 ), .C(FIFO_CLK_c), .D(n5677));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10851_4_lut (.I0(wr_addr_r[1]), .I1(wr_addr_r[4]), .I2(rp_sync_w[1]), 
            .I3(rp_sync_w[4]), .O(n12958));
    defparam i10851_4_lut.LUT_INIT = 16'hedb7;
    SB_DFF i272_273 (.Q(\REG.mem_2_14 ), .C(FIFO_CLK_c), .D(n5676));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14881_bdd_4_lut (.I0(n14881), .I1(n13853), .I2(n13852), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[30]));
    defparam n14881_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15571_bdd_4_lut (.I0(n15571), .I1(\REG.mem_5_13 ), .I2(\REG.mem_4_13 ), 
            .I3(rd_addr_r[1]), .O(n13884));
    defparam n15571_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10825_4_lut (.I0(wr_addr_r[3]), .I1(\wr_addr_r[0] ), .I2(rp_sync_w[3]), 
            .I3(rp_sync_w[0]), .O(n12932));
    defparam i10825_4_lut.LUT_INIT = 16'hedb7;
    SB_DFF i269_270 (.Q(\REG.mem_2_13 ), .C(FIFO_CLK_c), .D(n5675));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4574_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_14_2 ), .O(n6048));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4574_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12707 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_15 ), 
            .I2(\REG.mem_19_15 ), .I3(rd_addr_r[1]), .O(n14875));
    defparam rd_addr_r_0__bdd_4_lut_12707.LUT_INIT = 16'he4aa;
    SB_LUT4 n14875_bdd_4_lut (.I0(n14875), .I1(\REG.mem_17_15 ), .I2(\REG.mem_16_15 ), 
            .I3(rd_addr_r[1]), .O(n14878));
    defparam n14875_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13276 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_13 ), 
            .I2(\REG.mem_11_13 ), .I3(rd_addr_r[1]), .O(n15565));
    defparam rd_addr_r_0__bdd_4_lut_13276.LUT_INIT = 16'he4aa;
    SB_DFF i266_267 (.Q(\REG.mem_2_12 ), .C(FIFO_CLK_c), .D(n5674));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i263_264 (.Q(\REG.mem_2_11 ), .C(FIFO_CLK_c), .D(n5673));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i12230_3_lut (.I0(n12970), .I1(n12994), .I2(n8_adj_1377), 
            .I3(GND_net), .O(n14239));   // src/fifo_dc_32_lut_gen.v(300[45:114])
    defparam i12230_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 n15565_bdd_4_lut (.I0(n15565), .I1(\REG.mem_9_13 ), .I2(\REG.mem_8_13 ), 
            .I3(rd_addr_r[1]), .O(n13887));
    defparam n15565_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10939_4_lut (.I0(n12932), .I1(wr_addr_r[2]), .I2(n12958), 
            .I3(rp_sync_w[2]), .O(n13050));
    defparam i10939_4_lut.LUT_INIT = 16'hfefb;
    SB_LUT4 wr_addr_r_5__I_0_add_2_7_lut (.I0(n12209), .I1(\wr_addr_r[5] ), 
            .I2(n1_adj_1394[5]), .I3(n12106), .O(\afull_flag_impl.af_flag_nxt_w )) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_7_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 full_nxt_c_I_10_4_lut (.I0(n13050), .I1(n14239), .I2(wr_fifo_en_w), 
            .I3(dc32_fifo_full), .O(full_nxt_c_N_633));   // src/fifo_dc_32_lut_gen.v(300[45:114])
    defparam full_nxt_c_I_10_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12697 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_16 ), 
            .I2(\REG.mem_31_16 ), .I3(rd_addr_r[1]), .O(n14869));
    defparam rd_addr_r_0__bdd_4_lut_12697.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12488 (.I0(rd_addr_r[1]), .I1(n13312), 
            .I2(n13313), .I3(rd_addr_r[2]), .O(n14503));
    defparam rd_addr_r_1__bdd_4_lut_12488.LUT_INIT = 16'he4aa;
    SB_LUT4 n14503_bdd_4_lut (.I0(n14503), .I1(n13307), .I2(n13306), .I3(rd_addr_r[2]), 
            .O(n14506));
    defparam n14503_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12533 (.I0(rd_addr_r[3]), .I1(n14506), 
            .I2(n13058), .I3(rd_addr_r[4]), .O(n14539));
    defparam rd_addr_r_3__bdd_4_lut_12533.LUT_INIT = 16'he4aa;
    SB_LUT4 n14527_bdd_4_lut (.I0(n14527), .I1(n13812), .I2(n13650), .I3(rd_addr_r[3]), 
            .O(n14530));
    defparam n14527_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12400 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_4 ), 
            .I2(\REG.mem_19_4 ), .I3(rd_addr_r[1]), .O(n14497));
    defparam rd_addr_r_0__bdd_4_lut_12400.LUT_INIT = 16'he4aa;
    SB_LUT4 n14497_bdd_4_lut (.I0(n14497), .I1(\REG.mem_17_4 ), .I2(\REG.mem_16_4 ), 
            .I3(rd_addr_r[1]), .O(n14500));
    defparam n14497_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4110_2_lut_4_lut (.I0(rd_addr_r[0]), .I1(rd_addr_p1_w[0]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n5584));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4110_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 n14869_bdd_4_lut (.I0(n14869), .I1(\REG.mem_29_16 ), .I2(\REG.mem_28_16 ), 
            .I3(rd_addr_r[1]), .O(n14872));
    defparam n14869_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14539_bdd_4_lut (.I0(n14539), .I1(n13325), .I2(n13324), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[10]));
    defparam n14539_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4573_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_14_1 ), .O(n6047));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4573_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_13326 (.I0(rd_addr_r[3]), .I1(n15514), 
            .I2(n13706), .I3(rd_addr_r[4]), .O(n15553));
    defparam rd_addr_r_3__bdd_4_lut_13326.LUT_INIT = 16'he4aa;
    SB_LUT4 n15553_bdd_4_lut (.I0(n15553), .I1(n13691), .I2(n13690), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[26]));
    defparam n15553_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12692 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_19 ), 
            .I2(\REG.mem_11_19 ), .I3(rd_addr_r[1]), .O(n14863));
    defparam rd_addr_r_0__bdd_4_lut_12692.LUT_INIT = 16'he4aa;
    SB_DFF i260_261 (.Q(\REG.mem_2_10 ), .C(FIFO_CLK_c), .D(n5672));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i11307_3_lut (.I0(n15220), .I1(n15670), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13418));
    defparam i11307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_5__I_0_add_2_6_lut (.I0(n6_adj_1378), .I1(wr_addr_r[4]), 
            .I2(rp_sync_w[4]), .I3(n12105), .O(n8_adj_1373)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11252_3_lut (.I0(\REG.mem_24_22 ), .I1(\REG.mem_25_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13363));
    defparam i11252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_5__I_0_137_7_lut (.I0(GND_net), .I1(rd_grey_sync_r[5]), 
            .I2(GND_net), .I3(n12136), .O(rd_addr_p1_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11253_3_lut (.I0(\REG.mem_26_22 ), .I1(\REG.mem_27_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13364));
    defparam i11253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n14863_bdd_4_lut (.I0(n14863), .I1(\REG.mem_9_19 ), .I2(\REG.mem_8_19 ), 
            .I3(rd_addr_r[1]), .O(n13167));
    defparam n14863_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13271 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_6 ), 
            .I2(\REG.mem_3_6 ), .I3(rd_addr_r[1]), .O(n15547));
    defparam rd_addr_r_0__bdd_4_lut_13271.LUT_INIT = 16'he4aa;
    SB_DFF i257_258 (.Q(\REG.mem_2_9 ), .C(FIFO_CLK_c), .D(n5671));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i254_255 (.Q(\REG.mem_2_8 ), .C(FIFO_CLK_c), .D(n5670));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1265_1266 (.Q(\REG.mem_12_25 ), .C(FIFO_CLK_c), .D(n6007));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1262_1263 (.Q(\REG.mem_12_24 ), .C(FIFO_CLK_c), .D(n6006));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1259_1260 (.Q(\REG.mem_12_23 ), .C(FIFO_CLK_c), .D(n6005));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1256_1257 (.Q(\REG.mem_12_22 ), .C(FIFO_CLK_c), .D(n6004));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1253_1254 (.Q(\REG.mem_12_21 ), .C(FIFO_CLK_c), .D(n6003));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i251_252 (.Q(\REG.mem_2_7 ), .C(FIFO_CLK_c), .D(n5669));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12468 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_23 ), 
            .I2(\REG.mem_15_23 ), .I3(rd_addr_r[1]), .O(n14593));
    defparam rd_addr_r_0__bdd_4_lut_12468.LUT_INIT = 16'he4aa;
    SB_LUT4 i4572_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_14_0 ), .O(n6046));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4572_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11262_3_lut (.I0(\REG.mem_30_22 ), .I1(\REG.mem_31_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13373));
    defparam i11262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11261_3_lut (.I0(\REG.mem_28_22 ), .I1(\REG.mem_29_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13372));
    defparam i11261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11657_3_lut (.I0(\REG.mem_0_27 ), .I1(\REG.mem_1_27 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13768));
    defparam i11657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11658_3_lut (.I0(\REG.mem_2_27 ), .I1(\REG.mem_3_27 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13769));
    defparam i11658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12012_3_lut (.I0(\REG.mem_6_27 ), .I1(\REG.mem_7_27 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14123));
    defparam i12012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12011_3_lut (.I0(\REG.mem_4_27 ), .I1(\REG.mem_5_27 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14122));
    defparam i12011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n15547_bdd_4_lut (.I0(n15547), .I1(\REG.mem_1_6 ), .I2(\REG.mem_0_6 ), 
            .I3(rd_addr_r[1]), .O(n13890));
    defparam n15547_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12747 (.I0(rd_addr_r[1]), .I1(n13294), 
            .I2(n13295), .I3(rd_addr_r[2]), .O(n14857));
    defparam rd_addr_r_1__bdd_4_lut_12747.LUT_INIT = 16'he4aa;
    SB_LUT4 n14857_bdd_4_lut (.I0(n14857), .I1(n13289), .I2(n13288), .I3(rd_addr_r[2]), 
            .O(n13324));
    defparam n14857_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12702 (.I0(rd_addr_r[3]), .I1(n14848), 
            .I2(n13316), .I3(rd_addr_r[4]), .O(n14851));
    defparam rd_addr_r_3__bdd_4_lut_12702.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13256 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_21 ), 
            .I2(\REG.mem_15_21 ), .I3(rd_addr_r[1]), .O(n15541));
    defparam rd_addr_r_0__bdd_4_lut_13256.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_5__I_0_137_6_lut (.I0(GND_net), .I1(rd_addr_r[4]), 
            .I2(GND_net), .I3(n12135), .O(rd_addr_p1_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12062_3_lut (.I0(\REG.mem_16_27 ), .I1(\REG.mem_17_27 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14173));
    defparam i12062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12063_3_lut (.I0(\REG.mem_18_27 ), .I1(\REG.mem_19_27 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14174));
    defparam i12063_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rd_addr_r_5__I_0_137_6 (.CI(n12135), .I0(rd_addr_r[4]), .I1(GND_net), 
            .CO(n12136));
    SB_LUT4 rd_addr_r_5__I_0_137_5_lut (.I0(GND_net), .I1(rd_addr_r[3]), 
            .I2(GND_net), .I3(n12134), .O(rd_addr_p1_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rd_addr_r_5__I_0_137_5 (.CI(n12134), .I0(rd_addr_r[3]), .I1(GND_net), 
            .CO(n12135));
    SB_LUT4 rd_addr_r_5__I_0_137_4_lut (.I0(GND_net), .I1(rd_addr_r[2]), 
            .I2(GND_net), .I3(n12133), .O(rd_addr_p1_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_5__I_0_add_2_6 (.CI(n12105), .I0(wr_addr_r[4]), .I1(rp_sync_w[4]), 
            .CO(n12106));
    SB_LUT4 wr_addr_r_5__I_0_add_2_5_lut (.I0(wr_sig_diff0_w[2]), .I1(wr_addr_r[3]), 
            .I2(rp_sync_w[3]), .I3(n12104), .O(n7_adj_1372)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY wr_addr_r_5__I_0_add_2_5 (.CI(n12104), .I0(wr_addr_r[3]), .I1(rp_sync_w[3]), 
            .CO(n12105));
    SB_CARRY rd_addr_r_5__I_0_137_4 (.CI(n12133), .I0(rd_addr_r[2]), .I1(GND_net), 
            .CO(n12134));
    SB_LUT4 wr_addr_r_5__I_0_add_2_4_lut (.I0(GND_net), .I1(wr_addr_r[2]), 
            .I2(rp_sync_w[2]), .I3(n12103), .O(wr_sig_diff0_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_r_5__I_0_137_3_lut (.I0(GND_net), .I1(rd_addr_r[1]), 
            .I2(GND_net), .I3(n12132), .O(rd_addr_p1_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11237_3_lut (.I0(\REG.mem_8_2 ), .I1(\REG.mem_9_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13348));
    defparam i11237_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rd_addr_r_5__I_0_137_3 (.CI(n12132), .I0(rd_addr_r[1]), .I1(GND_net), 
            .CO(n12133));
    SB_LUT4 n14593_bdd_4_lut (.I0(n14593), .I1(\REG.mem_13_23 ), .I2(\REG.mem_12_23 ), 
            .I3(rd_addr_r[1]), .O(n14596));
    defparam n14593_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i248_249 (.Q(\REG.mem_2_6 ), .C(FIFO_CLK_c), .D(n5668));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14851_bdd_4_lut (.I0(n14851), .I1(n13304), .I2(n14842), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[7]));
    defparam n14851_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i245_246 (.Q(\REG.mem_2_5 ), .C(FIFO_CLK_c), .D(n5667));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i242_243 (.Q(\REG.mem_2_4 ), .C(FIFO_CLK_c), .D(n5666));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12387 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_12 ), 
            .I2(\REG.mem_23_12 ), .I3(rd_addr_r[1]), .O(n14491));
    defparam rd_addr_r_0__bdd_4_lut_12387.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_nxt_c_5__I_0_138_i1_2_lut_4_lut (.I0(rd_addr_r[0]), .I1(rd_addr_p1_w[0]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_5__N_573[1] ), .O(rd_grey_w[0]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_5__I_0_138_i1_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i11238_3_lut (.I0(\REG.mem_10_2 ), .I1(\REG.mem_11_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13349));
    defparam i11238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_nxt_c_5__I_0_136_i2_2_lut_4_lut (.I0(wr_addr_r[1]), .I1(wr_addr_p1_w[1]), 
            .I2(wr_fifo_en_w), .I3(\wr_addr_nxt_c[2] ), .O(wr_grey_w[1]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_5__I_0_136_i2_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i5457_2_lut_4_lut (.I0(wr_addr_r[1]), .I1(wr_addr_p1_w[1]), 
            .I2(wr_fifo_en_w), .I3(reset_per_frame), .O(n6931));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i5457_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 rd_addr_r_5__I_0_137_2_lut (.I0(GND_net), .I1(rd_addr_r[0]), 
            .I2(GND_net), .I3(VCC_net), .O(rd_addr_p1_w[0])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n15541_bdd_4_lut (.I0(n15541), .I1(\REG.mem_13_21 ), .I2(\REG.mem_12_21 ), 
            .I3(rd_addr_r[1]), .O(n15544));
    defparam n15541_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY rd_addr_r_5__I_0_137_2 (.CI(VCC_net), .I0(rd_addr_r[0]), .I1(GND_net), 
            .CO(n12132));
    SB_LUT4 wr_addr_r_5__I_0_128_7_lut (.I0(GND_net), .I1(\wr_addr_r[5] ), 
            .I2(GND_net), .I3(n12131), .O(wr_addr_p1_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_5__I_0_add_2_4 (.CI(n12103), .I0(wr_addr_r[2]), .I1(rp_sync_w[2]), 
            .CO(n12104));
    SB_LUT4 wr_addr_r_5__I_0_128_6_lut (.I0(GND_net), .I1(wr_addr_r[4]), 
            .I2(GND_net), .I3(n12130), .O(wr_addr_p1_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_5__I_0_128_6 (.CI(n12130), .I0(wr_addr_r[4]), .I1(GND_net), 
            .CO(n12131));
    SB_LUT4 wr_addr_r_5__I_0_128_5_lut (.I0(GND_net), .I1(wr_addr_r[3]), 
            .I2(GND_net), .I3(n12129), .O(wr_addr_p1_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11628_3_lut (.I0(\REG.mem_22_27 ), .I1(\REG.mem_23_27 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13739));
    defparam i11628_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY wr_addr_r_5__I_0_128_5 (.CI(n12129), .I0(wr_addr_r[3]), .I1(GND_net), 
            .CO(n12130));
    SB_LUT4 wr_addr_r_5__I_0_128_4_lut (.I0(GND_net), .I1(wr_addr_r[2]), 
            .I2(GND_net), .I3(n12128), .O(wr_addr_p1_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wr_addr_r_5__I_0_add_2_3_lut (.I0(n8993), .I1(wr_addr_r[1]), 
            .I2(rp_sync_w[1]), .I3(n12102), .O(n6_adj_1378)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY wr_addr_r_5__I_0_add_2_3 (.CI(n12102), .I0(wr_addr_r[1]), .I1(rp_sync_w[1]), 
            .CO(n12103));
    SB_CARRY wr_addr_r_5__I_0_128_4 (.CI(n12128), .I0(wr_addr_r[2]), .I1(GND_net), 
            .CO(n12129));
    SB_LUT4 wr_addr_r_5__I_0_add_2_2_lut (.I0(dc32_fifo_write_enable), .I1(\wr_addr_r[0] ), 
            .I2(rp_sync_w[0]), .I3(VCC_net), .O(n8993)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12682 (.I0(rd_addr_r[1]), .I1(n13897), 
            .I2(n13898), .I3(rd_addr_r[2]), .O(n14845));
    defparam rd_addr_r_1__bdd_4_lut_12682.LUT_INIT = 16'he4aa;
    SB_LUT4 i11627_3_lut (.I0(\REG.mem_20_27 ), .I1(\REG.mem_21_27 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13738));
    defparam i11627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n14845_bdd_4_lut (.I0(n14845), .I1(n13274), .I2(n13273), .I3(rd_addr_r[2]), 
            .O(n14848));
    defparam n14845_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13321 (.I0(rd_addr_r[1]), .I1(n13276), 
            .I2(n13277), .I3(rd_addr_r[2]), .O(n15535));
    defparam rd_addr_r_1__bdd_4_lut_13321.LUT_INIT = 16'he4aa;
    SB_LUT4 i4571_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_13_31 ), .O(n6045));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4571_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_addr_nxt_c_5__I_0_136_i1_2_lut_4_lut (.I0(wr_addr_r[1]), .I1(wr_addr_p1_w[1]), 
            .I2(wr_fifo_en_w), .I3(wr_addr_nxt_c[0]), .O(wr_grey_w[0]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_5__I_0_136_i1_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12672 (.I0(rd_addr_r[1]), .I1(n13240), 
            .I2(n13241), .I3(rd_addr_r[2]), .O(n14839));
    defparam rd_addr_r_1__bdd_4_lut_12672.LUT_INIT = 16'he4aa;
    SB_LUT4 n14839_bdd_4_lut (.I0(n14839), .I1(n13589), .I2(n13588), .I3(rd_addr_r[2]), 
            .O(n14842));
    defparam n14839_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_r_5__I_0_128_3_lut (.I0(GND_net), .I1(wr_addr_r[1]), 
            .I2(GND_net), .I3(n12127), .O(wr_addr_p1_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_5__I_0_add_2_2 (.CI(VCC_net), .I0(\wr_addr_r[0] ), 
            .I1(rp_sync_w[0]), .CO(n12102));
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_7_lut (.I0(rd_sig_diff0_w[3]), .I1(wp_sync2_r[5]), 
            .I2(n1[5]), .I3(n12070), .O(n6_adj_1379)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_7_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 n15535_bdd_4_lut (.I0(n15535), .I1(n13271), .I2(n13270), .I3(rd_addr_r[2]), 
            .O(n13892));
    defparam n15535_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13251 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_0 ), 
            .I2(\REG.mem_3_0 ), .I3(rd_addr_r[1]), .O(n15529));
    defparam rd_addr_r_0__bdd_4_lut_13251.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12677 (.I0(rd_addr_r[3]), .I1(n13891), 
            .I2(n13892), .I3(rd_addr_r[4]), .O(n14833));
    defparam rd_addr_r_3__bdd_4_lut_12677.LUT_INIT = 16'he4aa;
    SB_LUT4 n15529_bdd_4_lut (.I0(n15529), .I1(\REG.mem_1_0 ), .I2(\REG.mem_0_0 ), 
            .I3(rd_addr_r[1]), .O(n13425));
    defparam n15529_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY wr_addr_r_5__I_0_128_3 (.CI(n12127), .I0(wr_addr_r[1]), .I1(GND_net), 
            .CO(n12128));
    SB_LUT4 wr_addr_r_5__I_0_128_2_lut (.I0(GND_net), .I1(\wr_addr_r[0] ), 
            .I2(GND_net), .I3(VCC_net), .O(\wr_addr_p1_w[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4570_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_13_30 ), .O(n6044));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4570_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14833_bdd_4_lut (.I0(n14833), .I1(n13280), .I2(n14824), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[9]));
    defparam n14833_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_13306 (.I0(rd_addr_r[2]), .I1(n13827), 
            .I2(n13851), .I3(rd_addr_r[3]), .O(n15523));
    defparam rd_addr_r_2__bdd_4_lut_13306.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12662 (.I0(rd_addr_r[3]), .I1(n14818), 
            .I2(n13268), .I3(rd_addr_r[4]), .O(n14827));
    defparam rd_addr_r_3__bdd_4_lut_12662.LUT_INIT = 16'he4aa;
    SB_LUT4 n14827_bdd_4_lut (.I0(n14827), .I1(n13247), .I2(n14812), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[14]));
    defparam n14827_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12667 (.I0(rd_addr_r[1]), .I1(n13243), 
            .I2(n13244), .I3(rd_addr_r[2]), .O(n14821));
    defparam rd_addr_r_1__bdd_4_lut_12667.LUT_INIT = 16'he4aa;
    SB_LUT4 i4569_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_13_29 ), .O(n6043));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4569_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4568_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_13_28 ), .O(n6042));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4568_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15523_bdd_4_lut (.I0(n15523), .I1(n13662), .I2(n13794), .I3(rd_addr_r[3]), 
            .O(n15526));
    defparam n15523_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i239_240 (.Q(\REG.mem_2_3 ), .C(FIFO_CLK_c), .D(n5650));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4567_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_13_27 ), .O(n6041));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4567_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i65_66 (.Q(\REG.mem_0_9 ), .C(FIFO_CLK_c), .D(n5649));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i68_69 (.Q(\REG.mem_0_10 ), .C(FIFO_CLK_c), .D(n5642));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i71_72 (.Q(\REG.mem_0_11 ), .C(FIFO_CLK_c), .D(n5641));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1250_1251 (.Q(\REG.mem_12_20 ), .C(FIFO_CLK_c), .D(n6002));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13241 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_15 ), 
            .I2(\REG.mem_11_15 ), .I3(rd_addr_r[1]), .O(n15517));
    defparam rd_addr_r_0__bdd_4_lut_13241.LUT_INIT = 16'he4aa;
    SB_LUT4 n15517_bdd_4_lut (.I0(n15517), .I1(\REG.mem_9_15 ), .I2(\REG.mem_8_15 ), 
            .I3(rd_addr_r[1]), .O(n15520));
    defparam n15517_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14821_bdd_4_lut (.I0(n14821), .I1(n13238), .I2(n13237), .I3(rd_addr_r[2]), 
            .O(n14824));
    defparam n14821_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4148_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_0_24 ), .O(n5622));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4148_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4566_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_13_26 ), .O(n6040));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4566_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4565_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_13_25 ), .O(n6039));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4565_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1247_1248 (.Q(\REG.mem_12_19 ), .C(FIFO_CLK_c), .D(n6001));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1244_1245 (.Q(\REG.mem_12_18 ), .C(FIFO_CLK_c), .D(n6000));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1241_1242 (.Q(\REG.mem_12_17 ), .C(FIFO_CLK_c), .D(n5999));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1238_1239 (.Q(\REG.mem_12_16 ), .C(FIFO_CLK_c), .D(n5998));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i236_237 (.Q(\REG.mem_2_2 ), .C(FIFO_CLK_c), .D(n5640));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12652 (.I0(rd_addr_r[1]), .I1(n13228), 
            .I2(n13229), .I3(rd_addr_r[2]), .O(n14815));
    defparam rd_addr_r_1__bdd_4_lut_12652.LUT_INIT = 16'he4aa;
    SB_LUT4 n14815_bdd_4_lut (.I0(n14815), .I1(n13226), .I2(n13225), .I3(rd_addr_r[2]), 
            .O(n14818));
    defparam n14815_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13246 (.I0(rd_addr_r[1]), .I1(n13633), 
            .I2(n13634), .I3(rd_addr_r[2]), .O(n15511));
    defparam rd_addr_r_1__bdd_4_lut_13246.LUT_INIT = 16'he4aa;
    SB_LUT4 i4564_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_13_24 ), .O(n6038));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4564_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12647 (.I0(rd_addr_r[1]), .I1(n13216), 
            .I2(n13217), .I3(rd_addr_r[2]), .O(n14809));
    defparam rd_addr_r_1__bdd_4_lut_12647.LUT_INIT = 16'he4aa;
    SB_LUT4 n15511_bdd_4_lut (.I0(n15511), .I1(n13712), .I2(n13711), .I3(rd_addr_r[2]), 
            .O(n15514));
    defparam n15511_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14809_bdd_4_lut (.I0(n14809), .I1(n13214), .I2(n13213), .I3(rd_addr_r[2]), 
            .O(n14812));
    defparam n14809_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11285_3_lut (.I0(\REG.mem_16_1 ), .I1(\REG.mem_17_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13396));
    defparam i11285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11286_3_lut (.I0(\REG.mem_18_1 ), .I1(\REG.mem_19_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13397));
    defparam i11286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12657 (.I0(rd_addr_r[3]), .I1(n13963), 
            .I2(n13964), .I3(rd_addr_r[4]), .O(n14803));
    defparam rd_addr_r_3__bdd_4_lut_12657.LUT_INIT = 16'he4aa;
    SB_LUT4 i4095_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_0_2 ), .O(n5569));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4095_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14803_bdd_4_lut (.I0(n14803), .I1(n13211), .I2(n13210), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[18]));
    defparam n14803_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12642 (.I0(rd_addr_r[1]), .I1(n13546), 
            .I2(n13547), .I3(rd_addr_r[2]), .O(n14797));
    defparam rd_addr_r_1__bdd_4_lut_12642.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13226 (.I0(rd_addr_r[1]), .I1(n13747), 
            .I2(n13748), .I3(rd_addr_r[2]), .O(n15505));
    defparam rd_addr_r_1__bdd_4_lut_13226.LUT_INIT = 16'he4aa;
    SB_LUT4 n15505_bdd_4_lut (.I0(n15505), .I1(n14135), .I2(n14134), .I3(rd_addr_r[2]), 
            .O(n13433));
    defparam n15505_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14797_bdd_4_lut (.I0(n14797), .I1(n14162), .I2(n14161), .I3(rd_addr_r[2]), 
            .O(n14800));
    defparam n14797_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4563_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_13_23 ), .O(n6037));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4563_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4562_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_13_22 ), .O(n6036));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4562_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i74_75 (.Q(\REG.mem_0_12 ), .C(FIFO_CLK_c), .D(n5639));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i77_78 (.Q(\REG.mem_0_13 ), .C(FIFO_CLK_c), .D(n5638));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i80_81 (.Q(\REG.mem_0_14 ), .C(FIFO_CLK_c), .D(n5637));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i83_84 (.Q(\REG.mem_0_15 ), .C(FIFO_CLK_c), .D(n5634));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i86_87 (.Q(\REG.mem_0_16 ), .C(FIFO_CLK_c), .D(n5633));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i89_90 (.Q(\REG.mem_0_17 ), .C(FIFO_CLK_c), .D(n5632));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i59_60 (.Q(\REG.mem_0_7 ), .C(FIFO_CLK_c), .D(n5631));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i92_93 (.Q(\REG.mem_0_18 ), .C(FIFO_CLK_c), .D(n5630));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i95_96 (.Q(\REG.mem_0_19 ), .C(FIFO_CLK_c), .D(n5629));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13221 (.I0(rd_addr_r[1]), .I1(n13336), 
            .I2(n13337), .I3(rd_addr_r[2]), .O(n15493));
    defparam rd_addr_r_1__bdd_4_lut_13221.LUT_INIT = 16'he4aa;
    SB_LUT4 n15493_bdd_4_lut (.I0(n15493), .I1(n13844), .I2(n13843), .I3(rd_addr_r[2]), 
            .O(n15496));
    defparam n15493_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13231 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_13 ), 
            .I2(\REG.mem_15_13 ), .I3(rd_addr_r[1]), .O(n15487));
    defparam rd_addr_r_0__bdd_4_lut_13231.LUT_INIT = 16'he4aa;
    SB_LUT4 n15487_bdd_4_lut (.I0(n15487), .I1(\REG.mem_13_13 ), .I2(\REG.mem_12_13 ), 
            .I3(rd_addr_r[1]), .O(n13902));
    defparam n15487_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12632 (.I0(rd_addr_r[1]), .I1(n13108), 
            .I2(n13109), .I3(rd_addr_r[2]), .O(n14791));
    defparam rd_addr_r_1__bdd_4_lut_12632.LUT_INIT = 16'he4aa;
    SB_LUT4 n14791_bdd_4_lut (.I0(n14791), .I1(n13097), .I2(n13096), .I3(rd_addr_r[2]), 
            .O(n14794));
    defparam n14791_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i98_99 (.Q(\REG.mem_0_20 ), .C(FIFO_CLK_c), .D(n5628));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4561_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_13_21 ), .O(n6035));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4561_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12687 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_0 ), 
            .I2(\REG.mem_27_0 ), .I3(rd_addr_r[1]), .O(n14785));
    defparam rd_addr_r_0__bdd_4_lut_12687.LUT_INIT = 16'he4aa;
    SB_DFFE \REG.out_raw_i0_i2  (.Q(\dc32_fifo_data_out[1] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[1]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_LUT4 n14785_bdd_4_lut (.I0(n14785), .I1(\REG.mem_25_0 ), .I2(\REG.mem_24_0 ), 
            .I3(rd_addr_r[1]), .O(n14788));
    defparam n14785_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13206 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_16 ), 
            .I2(\REG.mem_19_16 ), .I3(rd_addr_r[1]), .O(n15481));
    defparam rd_addr_r_0__bdd_4_lut_13206.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12622 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_11 ), 
            .I2(\REG.mem_11_11 ), .I3(rd_addr_r[1]), .O(n14779));
    defparam rd_addr_r_0__bdd_4_lut_12622.LUT_INIT = 16'he4aa;
    SB_LUT4 n14779_bdd_4_lut (.I0(n14779), .I1(\REG.mem_9_11 ), .I2(\REG.mem_8_11 ), 
            .I3(rd_addr_r[1]), .O(n14782));
    defparam n14779_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15481_bdd_4_lut (.I0(n15481), .I1(\REG.mem_17_16 ), .I2(\REG.mem_16_16 ), 
            .I3(rd_addr_r[1]), .O(n15484));
    defparam n15481_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \REG.out_raw_i0_i3  (.Q(\dc32_fifo_data_out[2] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[2]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i4  (.Q(\dc32_fifo_data_out[3] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[3]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i5  (.Q(\dc32_fifo_data_out[4] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[4]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i6  (.Q(\dc32_fifo_data_out[5] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[5]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i7  (.Q(\dc32_fifo_data_out[6] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[6]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i8  (.Q(\dc32_fifo_data_out[7] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[7]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i9  (.Q(\dc32_fifo_data_out[8] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[8]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i10  (.Q(\dc32_fifo_data_out[9] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[9]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i11  (.Q(\dc32_fifo_data_out[10] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[10]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i12  (.Q(\dc32_fifo_data_out[11] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[11]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i13  (.Q(\dc32_fifo_data_out[12] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[12]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i14  (.Q(\dc32_fifo_data_out[13] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[13]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i15  (.Q(\dc32_fifo_data_out[14] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[14]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i16  (.Q(\dc32_fifo_data_out[15] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[15]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i17  (.Q(\dc32_fifo_data_out[16] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[16]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i18  (.Q(\dc32_fifo_data_out[17] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[17]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i19  (.Q(\dc32_fifo_data_out[18] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[18]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i20  (.Q(\dc32_fifo_data_out[19] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[19]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i21  (.Q(\dc32_fifo_data_out[20] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[20]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i22  (.Q(\dc32_fifo_data_out[21] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[21]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i23  (.Q(\dc32_fifo_data_out[22] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[22]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i24  (.Q(\dc32_fifo_data_out[23] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[23]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i25  (.Q(\dc32_fifo_data_out[24] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[24]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i26  (.Q(\dc32_fifo_data_out[25] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[25]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i27  (.Q(\dc32_fifo_data_out[26] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[26]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i28  (.Q(\dc32_fifo_data_out[27] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[27]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i29  (.Q(\dc32_fifo_data_out[28] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[28]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i30  (.Q(\dc32_fifo_data_out[29] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[29]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i31  (.Q(\dc32_fifo_data_out[30] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[30]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i32  (.Q(\dc32_fifo_data_out[31] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[31]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFF i1235_1236 (.Q(\REG.mem_12_15 ), .C(FIFO_CLK_c), .D(n5997));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4560_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_13_20 ), .O(n6034));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4560_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12617 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_19 ), 
            .I2(\REG.mem_15_19 ), .I3(rd_addr_r[1]), .O(n14773));
    defparam rd_addr_r_0__bdd_4_lut_12617.LUT_INIT = 16'he4aa;
    SB_LUT4 n14773_bdd_4_lut (.I0(n14773), .I1(\REG.mem_13_19 ), .I2(\REG.mem_12_19 ), 
            .I3(rd_addr_r[1]), .O(n13170));
    defparam n14773_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_6_lut (.I0(n46), .I1(wp_sync_w[4]), 
            .I2(n1[4]), .I3(n12069), .O(n7_adj_3)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_6_lut.LUT_INIT = 16'hebbe;
    SB_CARRY wp_sync2_r_5__I_0_135_add_2_6 (.CI(n12069), .I0(wp_sync_w[4]), 
            .I1(n1[4]), .CO(n12070));
    SB_CARRY wr_addr_r_5__I_0_128_2 (.CI(VCC_net), .I0(\wr_addr_r[0] ), 
            .I1(GND_net), .CO(n12127));
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_5_lut (.I0(GND_net), .I1(wp_sync_w[3]), 
            .I2(n1[3]), .I3(n12068), .O(rd_sig_diff0_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wp_sync2_r_5__I_0_135_add_2_5 (.CI(n12068), .I0(wp_sync_w[3]), 
            .I1(n1[3]), .CO(n12069));
    SB_DFF i1232_1233 (.Q(\REG.mem_12_14 ), .C(FIFO_CLK_c), .D(n5996));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_4_lut (.I0(n6_adj_1379), .I1(wp_sync_w[2]), 
            .I2(n1[2]), .I3(n12067), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 EnabledDecoder_2_i21_2_lut (.I0(n13_c), .I1(wr_addr_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i21_2_lut.LUT_INIT = 16'h2222;
    SB_DFF i1229_1230 (.Q(\REG.mem_12_13 ), .C(FIFO_CLK_c), .D(n5995));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1226_1227 (.Q(\REG.mem_12_12 ), .C(FIFO_CLK_c), .D(n5994));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1223_1224 (.Q(\REG.mem_12_11 ), .C(FIFO_CLK_c), .D(n5993));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1220_1221 (.Q(\REG.mem_12_10 ), .C(FIFO_CLK_c), .D(n5992));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i233_234 (.Q(\REG.mem_2_1 ), .C(FIFO_CLK_c), .D(n5627));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4559_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_13_19 ), .O(n6033));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4559_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY wp_sync2_r_5__I_0_135_add_2_4 (.CI(n12067), .I0(wp_sync_w[2]), 
            .I1(n1[2]), .CO(n12068));
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_3_lut (.I0(n49), .I1(wp_sync_w[1]), 
            .I2(n1[1]), .I3(n12066), .O(n46)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY wp_sync2_r_5__I_0_135_add_2_3 (.CI(n12066), .I0(wp_sync_w[1]), 
            .I1(n1[1]), .CO(n12067));
    SB_DFF i230_231 (.Q(\REG.mem_2_0 ), .C(FIFO_CLK_c), .D(n5626));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1217_1218 (.Q(\REG.mem_12_9 ), .C(FIFO_CLK_c), .D(n5991));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1214_1215 (.Q(\REG.mem_12_8 ), .C(FIFO_CLK_c), .D(n5990));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1211_1212 (.Q(\REG.mem_12_7 ), .C(FIFO_CLK_c), .D(n5989));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_2_lut (.I0(n25), .I1(wp_sync_w[0]), 
            .I2(n1[0]), .I3(VCC_net), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12612 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_5 ), 
            .I2(\REG.mem_27_5 ), .I3(rd_addr_r[1]), .O(n14767));
    defparam rd_addr_r_0__bdd_4_lut_12612.LUT_INIT = 16'he4aa;
    SB_LUT4 n14767_bdd_4_lut (.I0(n14767), .I1(\REG.mem_25_5 ), .I2(\REG.mem_24_5 ), 
            .I3(rd_addr_r[1]), .O(n14770));
    defparam n14767_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1208_1209 (.Q(\REG.mem_12_6 ), .C(FIFO_CLK_c), .D(n5988));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i11292_3_lut (.I0(\REG.mem_22_1 ), .I1(\REG.mem_23_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13403));
    defparam i11292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13211 (.I0(rd_addr_r[1]), .I1(n13735), 
            .I2(n13736), .I3(rd_addr_r[2]), .O(n15469));
    defparam rd_addr_r_1__bdd_4_lut_13211.LUT_INIT = 16'he4aa;
    SB_LUT4 i11291_3_lut (.I0(\REG.mem_20_1 ), .I1(\REG.mem_21_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13402));
    defparam i11291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12607 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_19 ), 
            .I2(\REG.mem_19_19 ), .I3(rd_addr_r[1]), .O(n14761));
    defparam rd_addr_r_0__bdd_4_lut_12607.LUT_INIT = 16'he4aa;
    SB_LUT4 n14761_bdd_4_lut (.I0(n14761), .I1(\REG.mem_17_19 ), .I2(\REG.mem_16_19 ), 
            .I3(rd_addr_r[1]), .O(n14764));
    defparam n14761_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11247_3_lut (.I0(\REG.mem_14_2 ), .I1(\REG.mem_15_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13358));
    defparam i11247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12602 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_5 ), 
            .I2(\REG.mem_31_5 ), .I3(rd_addr_r[1]), .O(n14755));
    defparam rd_addr_r_0__bdd_4_lut_12602.LUT_INIT = 16'he4aa;
    SB_LUT4 i11246_3_lut (.I0(\REG.mem_12_2 ), .I1(\REG.mem_13_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13357));
    defparam i11246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n15469_bdd_4_lut (.I0(n15469), .I1(n14180), .I2(n14179), .I3(rd_addr_r[2]), 
            .O(n15472));
    defparam n15469_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14755_bdd_4_lut (.I0(n14755), .I1(\REG.mem_29_5 ), .I2(\REG.mem_28_5 ), 
            .I3(rd_addr_r[1]), .O(n14758));
    defparam n14755_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i101_102 (.Q(\REG.mem_0_21 ), .C(FIFO_CLK_c), .D(n5625));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1205_1206 (.Q(\REG.mem_12_5 ), .C(FIFO_CLK_c), .D(n5987));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13201 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_8 ), 
            .I2(\REG.mem_15_8 ), .I3(rd_addr_r[1]), .O(n15463));
    defparam rd_addr_r_0__bdd_4_lut_13201.LUT_INIT = 16'he4aa;
    SB_DFF i1202_1203 (.Q(\REG.mem_12_4 ), .C(FIFO_CLK_c), .D(n5986));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1199_1200 (.Q(\REG.mem_12_3 ), .C(FIFO_CLK_c), .D(n5985));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1196_1197 (.Q(\REG.mem_12_2 ), .C(FIFO_CLK_c), .D(n5984));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1193_1194 (.Q(\REG.mem_12_1 ), .C(FIFO_CLK_c), .D(n5983));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1190_1191 (.Q(\REG.mem_12_0 ), .C(FIFO_CLK_c), .D(n5982));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i104_105 (.Q(\REG.mem_0_22 ), .C(FIFO_CLK_c), .D(n5624));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12597 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_0 ), 
            .I2(\REG.mem_31_0 ), .I3(rd_addr_r[1]), .O(n14749));
    defparam rd_addr_r_0__bdd_4_lut_12597.LUT_INIT = 16'he4aa;
    SB_DFF i107_108 (.Q(\REG.mem_0_23 ), .C(FIFO_CLK_c), .D(n5623));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n15463_bdd_4_lut (.I0(n15463), .I1(\REG.mem_13_8 ), .I2(\REG.mem_12_8 ), 
            .I3(rd_addr_r[1]), .O(n15466));
    defparam n15463_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14749_bdd_4_lut (.I0(n14749), .I1(\REG.mem_29_0 ), .I2(\REG.mem_28_0 ), 
            .I3(rd_addr_r[1]), .O(n14752));
    defparam n14749_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i110_111 (.Q(\REG.mem_0_24 ), .C(FIFO_CLK_c), .D(n5622));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i113_114 (.Q(\REG.mem_0_25 ), .C(FIFO_CLK_c), .D(n5621));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i116_117 (.Q(\REG.mem_0_26 ), .C(FIFO_CLK_c), .D(n5620));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1187_1188 (.Q(\REG.mem_11_31 ), .C(FIFO_CLK_c), .D(n5981));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12627 (.I0(rd_addr_r[1]), .I1(n14137), 
            .I2(n14138), .I3(rd_addr_r[2]), .O(n14743));
    defparam rd_addr_r_1__bdd_4_lut_12627.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13191 (.I0(rd_addr_r[1]), .I1(n14155), 
            .I2(n14156), .I3(rd_addr_r[2]), .O(n15457));
    defparam rd_addr_r_1__bdd_4_lut_13191.LUT_INIT = 16'he4aa;
    SB_LUT4 n14743_bdd_4_lut (.I0(n14743), .I1(n14132), .I2(n14131), .I3(rd_addr_r[2]), 
            .O(n14746));
    defparam n14743_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4558_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_13_18 ), .O(n6032));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4558_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15457_bdd_4_lut (.I0(n15457), .I1(n14144), .I2(n14143), .I3(rd_addr_r[2]), 
            .O(n13139));
    defparam n15457_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4557_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_13_17 ), .O(n6031));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4557_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4556_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_13_16 ), .O(n6030));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4556_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12592 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_23 ), 
            .I2(\REG.mem_3_23 ), .I3(rd_addr_r[1]), .O(n14725));
    defparam rd_addr_r_0__bdd_4_lut_12592.LUT_INIT = 16'he4aa;
    SB_LUT4 n14725_bdd_4_lut (.I0(n14725), .I1(\REG.mem_1_23 ), .I2(\REG.mem_0_23 ), 
            .I3(rd_addr_r[1]), .O(n14728));
    defparam n14725_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4555_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_13_15 ), .O(n6029));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4555_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1184_1185 (.Q(\REG.mem_11_30 ), .C(FIFO_CLK_c), .D(n5980));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14533_bdd_4_lut (.I0(n14533), .I1(\REG.mem_17_23 ), .I2(\REG.mem_16_23 ), 
            .I3(rd_addr_r[1]), .O(n14536));
    defparam n14533_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12573 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_19 ), 
            .I2(\REG.mem_23_19 ), .I3(rd_addr_r[1]), .O(n14719));
    defparam rd_addr_r_0__bdd_4_lut_12573.LUT_INIT = 16'he4aa;
    SB_LUT4 n14719_bdd_4_lut (.I0(n14719), .I1(\REG.mem_21_19 ), .I2(\REG.mem_20_19 ), 
            .I3(rd_addr_r[1]), .O(n14722));
    defparam n14719_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13186 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_6 ), 
            .I2(\REG.mem_7_6 ), .I3(rd_addr_r[1]), .O(n15445));
    defparam rd_addr_r_0__bdd_4_lut_13186.LUT_INIT = 16'he4aa;
    SB_LUT4 n15445_bdd_4_lut (.I0(n15445), .I1(\REG.mem_5_6 ), .I2(\REG.mem_4_6 ), 
            .I3(rd_addr_r[1]), .O(n13911));
    defparam n15445_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1181_1182 (.Q(\REG.mem_11_29 ), .C(FIFO_CLK_c), .D(n5979));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12568 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_29 ), 
            .I2(\REG.mem_11_29 ), .I3(rd_addr_r[1]), .O(n14713));
    defparam rd_addr_r_0__bdd_4_lut_12568.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12433 (.I0(rd_addr_r[2]), .I1(n13767), 
            .I2(n13830), .I3(rd_addr_r[3]), .O(n14527));
    defparam rd_addr_r_2__bdd_4_lut_12433.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13171 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_13 ), 
            .I2(\REG.mem_23_13 ), .I3(rd_addr_r[1]), .O(n15439));
    defparam rd_addr_r_0__bdd_4_lut_13171.LUT_INIT = 16'he4aa;
    SB_DFF i1178_1179 (.Q(\REG.mem_11_28 ), .C(FIFO_CLK_c), .D(n5978));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1175_1176 (.Q(\REG.mem_11_27 ), .C(FIFO_CLK_c), .D(n5977));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1172_1173 (.Q(\REG.mem_11_26 ), .C(FIFO_CLK_c), .D(n5976));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1169_1170 (.Q(\REG.mem_11_25 ), .C(FIFO_CLK_c), .D(n5975));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1166_1167 (.Q(\REG.mem_11_24 ), .C(FIFO_CLK_c), .D(n5974));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n15439_bdd_4_lut (.I0(n15439), .I1(\REG.mem_21_13 ), .I2(\REG.mem_20_13 ), 
            .I3(rd_addr_r[1]), .O(n13914));
    defparam n15439_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14713_bdd_4_lut (.I0(n14713), .I1(\REG.mem_9_29 ), .I2(\REG.mem_8_29 ), 
            .I3(rd_addr_r[1]), .O(n14716));
    defparam n14713_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1163_1164 (.Q(\REG.mem_11_23 ), .C(FIFO_CLK_c), .D(n5973));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12732 (.I0(rd_addr_r[2]), .I1(n13974), 
            .I2(n13998), .I3(rd_addr_r[3]), .O(n14707));
    defparam rd_addr_r_2__bdd_4_lut_12732.LUT_INIT = 16'he4aa;
    SB_LUT4 n14707_bdd_4_lut (.I0(n14707), .I1(n13632), .I2(n13926), .I3(rd_addr_r[3]), 
            .O(n14710));
    defparam n14707_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4554_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_13_14 ), .O(n6028));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4554_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1160_1161 (.Q(\REG.mem_11_22 ), .C(FIFO_CLK_c), .D(n5972));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12563 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_19 ), 
            .I2(\REG.mem_27_19 ), .I3(rd_addr_r[1]), .O(n14701));
    defparam rd_addr_r_0__bdd_4_lut_12563.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13166 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_13 ), 
            .I2(\REG.mem_27_13 ), .I3(rd_addr_r[1]), .O(n15427));
    defparam rd_addr_r_0__bdd_4_lut_13166.LUT_INIT = 16'he4aa;
    SB_LUT4 n14701_bdd_4_lut (.I0(n14701), .I1(\REG.mem_25_19 ), .I2(\REG.mem_24_19 ), 
            .I3(rd_addr_r[1]), .O(n14704));
    defparam n14701_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15427_bdd_4_lut (.I0(n15427), .I1(\REG.mem_25_13 ), .I2(\REG.mem_24_13 ), 
            .I3(rd_addr_r[1]), .O(n13917));
    defparam n15427_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i45_2_lut_3_lut (.I0(n12_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n29));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i45_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i11583_3_lut (.I0(n14716), .I1(n15748), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13694));
    defparam i11583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13156 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_28 ), 
            .I2(\REG.mem_19_28 ), .I3(rd_addr_r[1]), .O(n15421));
    defparam rd_addr_r_0__bdd_4_lut_13156.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12558 (.I0(rd_addr_r[2]), .I1(n13980), 
            .I2(n14004), .I3(rd_addr_r[3]), .O(n14695));
    defparam rd_addr_r_2__bdd_4_lut_12558.LUT_INIT = 16'he4aa;
    SB_LUT4 i4553_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_13_13 ), .O(n6027));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4553_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11618_3_lut (.I0(n14632), .I1(n15778), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13729));
    defparam i11618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut (.I0(rd_addr_r[0]), .I1(\REG.mem_22_4 ), 
            .I2(\REG.mem_23_4 ), .I3(rd_addr_r[1]), .O(n16225));
    defparam rd_addr_r_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n16225_bdd_4_lut (.I0(n16225), .I1(\REG.mem_21_4 ), .I2(\REG.mem_20_4 ), 
            .I3(rd_addr_r[1]), .O(n16228));
    defparam n16225_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4552_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_13_12 ), .O(n6026));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4552_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11210_3_lut (.I0(\REG.mem_8_17 ), .I1(\REG.mem_9_17 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13321));
    defparam i11210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n15421_bdd_4_lut (.I0(n15421), .I1(\REG.mem_17_28 ), .I2(\REG.mem_16_28 ), 
            .I3(rd_addr_r[1]), .O(n13920));
    defparam n15421_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut (.I0(rd_addr_r[2]), .I1(n15094), .I2(n14872), 
            .I3(rd_addr_r[3]), .O(n16219));
    defparam rd_addr_r_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n14695_bdd_4_lut (.I0(n14695), .I1(n13947), .I2(n13920), .I3(rd_addr_r[3]), 
            .O(n14698));
    defparam n14695_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16219_bdd_4_lut (.I0(n16219), .I1(n15274), .I2(n15484), .I3(rd_addr_r[3]), 
            .O(n16222));
    defparam n16219_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11211_3_lut (.I0(\REG.mem_10_17 ), .I1(\REG.mem_11_17 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13322));
    defparam i11211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11325_3_lut (.I0(n16060), .I1(n15244), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13436));
    defparam i11325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10950_3_lut (.I0(\REG.mem_14_17 ), .I1(\REG.mem_15_17 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13061));
    defparam i10950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13151 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_24 ), 
            .I2(\REG.mem_3_24 ), .I3(rd_addr_r[1]), .O(n15415));
    defparam rd_addr_r_0__bdd_4_lut_13151.LUT_INIT = 16'he4aa;
    SB_LUT4 i10949_3_lut (.I0(\REG.mem_12_17 ), .I1(\REG.mem_13_17 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13060));
    defparam i10949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12553 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_19 ), 
            .I2(\REG.mem_31_19 ), .I3(rd_addr_r[1]), .O(n14689));
    defparam rd_addr_r_0__bdd_4_lut_12553.LUT_INIT = 16'he4aa;
    SB_LUT4 n14689_bdd_4_lut (.I0(n14689), .I1(\REG.mem_29_19 ), .I2(\REG.mem_28_19 ), 
            .I3(rd_addr_r[1]), .O(n14692));
    defparam n14689_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13820 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_23 ), 
            .I2(\REG.mem_23_23 ), .I3(rd_addr_r[1]), .O(n16213));
    defparam rd_addr_r_0__bdd_4_lut_13820.LUT_INIT = 16'he4aa;
    SB_LUT4 i4551_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_13_11 ), .O(n6025));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4551_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15415_bdd_4_lut (.I0(n15415), .I1(\REG.mem_1_24 ), .I2(\REG.mem_0_24 ), 
            .I3(rd_addr_r[1]), .O(n13923));
    defparam n15415_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16213_bdd_4_lut (.I0(n16213), .I1(\REG.mem_21_23 ), .I2(\REG.mem_20_23 ), 
            .I3(rd_addr_r[1]), .O(n16216));
    defparam n16213_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10973_3_lut (.I0(\REG.mem_16_17 ), .I1(\REG.mem_17_17 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13084));
    defparam i10973_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1157_1158 (.Q(\REG.mem_11_21 ), .C(FIFO_CLK_c), .D(n5971));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4550_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_13_10 ), .O(n6024));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4550_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4549_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_13_9 ), .O(n6023));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4549_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1154_1155 (.Q(\REG.mem_11_20 ), .C(FIFO_CLK_c), .D(n5970));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13810 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_31 ), 
            .I2(\REG.mem_7_31 ), .I3(rd_addr_r[1]), .O(n16207));
    defparam rd_addr_r_0__bdd_4_lut_13810.LUT_INIT = 16'he4aa;
    SB_LUT4 n16207_bdd_4_lut (.I0(n16207), .I1(\REG.mem_5_31 ), .I2(\REG.mem_4_31 ), 
            .I3(rd_addr_r[1]), .O(n16210));
    defparam n16207_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12548 (.I0(rd_addr_r[2]), .I1(n14016), 
            .I2(n14025), .I3(rd_addr_r[3]), .O(n14683));
    defparam rd_addr_r_2__bdd_4_lut_12548.LUT_INIT = 16'he4aa;
    SB_DFF i119_120 (.Q(\REG.mem_0_27 ), .C(FIFO_CLK_c), .D(n5617));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10974_3_lut (.I0(\REG.mem_18_17 ), .I1(\REG.mem_19_17 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13085));
    defparam i10974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13146 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_15 ), 
            .I2(\REG.mem_15_15 ), .I3(rd_addr_r[1]), .O(n15403));
    defparam rd_addr_r_0__bdd_4_lut_13146.LUT_INIT = 16'he4aa;
    SB_LUT4 i4548_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_13_8 ), .O(n6022));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4548_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14683_bdd_4_lut (.I0(n14683), .I1(n14013), .I2(n14007), .I3(rd_addr_r[3]), 
            .O(n14686));
    defparam n14683_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12637 (.I0(rd_addr_r[3]), .I1(n14662), 
            .I2(n13124), .I3(rd_addr_r[4]), .O(n14677));
    defparam rd_addr_r_3__bdd_4_lut_12637.LUT_INIT = 16'he4aa;
    SB_LUT4 n14677_bdd_4_lut (.I0(n14677), .I1(n13121), .I2(n14650), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[11]));
    defparam n14677_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15403_bdd_4_lut (.I0(n15403), .I1(\REG.mem_13_15 ), .I2(\REG.mem_12_15 ), 
            .I3(rd_addr_r[1]), .O(n15406));
    defparam n15403_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i122_123 (.Q(\REG.mem_0_28 ), .C(FIFO_CLK_c), .D(n5616));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i125_126 (.Q(\REG.mem_0_29 ), .C(FIFO_CLK_c), .D(n5614));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFSR rd_grey_sync_r__i1 (.Q(rd_grey_sync_r[1]), .C(SLM_CLK_c), .D(rd_grey_w[1]), 
            .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i2 (.Q(rd_grey_sync_r[2]), .C(SLM_CLK_c), .D(rd_grey_w[2]), 
            .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i3 (.Q(rd_grey_sync_r[3]), .C(SLM_CLK_c), .D(rd_grey_w[3]), 
            .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i4 (.Q(rd_grey_sync_r[4]), .C(SLM_CLK_c), .D(rd_grey_w[4]), 
            .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR wr_grey_sync_r__i1 (.Q(\wr_grey_sync_r[1] ), .C(FIFO_CLK_c), 
            .D(wr_grey_w[1]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_LUT4 EnabledDecoder_2_i55_2_lut_3_lut (.I0(n15), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n24));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i55_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13805 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_31 ), 
            .I2(\REG.mem_19_31 ), .I3(rd_addr_r[1]), .O(n16195));
    defparam rd_addr_r_0__bdd_4_lut_13805.LUT_INIT = 16'he4aa;
    SB_LUT4 n16195_bdd_4_lut (.I0(n16195), .I1(\REG.mem_17_31 ), .I2(\REG.mem_16_31 ), 
            .I3(rd_addr_r[1]), .O(n16198));
    defparam n16195_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12538 (.I0(rd_addr_r[2]), .I1(n13464), 
            .I2(n13479), .I3(rd_addr_r[3]), .O(n14671));
    defparam rd_addr_r_2__bdd_4_lut_12538.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i44_2_lut_3_lut (.I0(n12_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n13));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i44_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13136 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_8 ), 
            .I2(\REG.mem_19_8 ), .I3(rd_addr_r[1]), .O(n15397));
    defparam rd_addr_r_0__bdd_4_lut_13136.LUT_INIT = 16'he4aa;
    SB_LUT4 n15397_bdd_4_lut (.I0(n15397), .I1(\REG.mem_17_8 ), .I2(\REG.mem_16_8 ), 
            .I3(rd_addr_r[1]), .O(n13926));
    defparam n15397_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12463 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_18 ), 
            .I2(\REG.mem_3_18 ), .I3(rd_addr_r[1]), .O(n14581));
    defparam rd_addr_r_0__bdd_4_lut_12463.LUT_INIT = 16'he4aa;
    SB_LUT4 i4547_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_13_7 ), .O(n6021));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4547_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i54_2_lut_3_lut (.I0(n15), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n8_adj_4));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i54_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 n14671_bdd_4_lut (.I0(n14671), .I1(n13452), .I2(n13425), .I3(rd_addr_r[3]), 
            .O(n14674));
    defparam n14671_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4175_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_0_9 ), .O(n5649));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4175_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13795 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_31 ), 
            .I2(\REG.mem_23_31 ), .I3(rd_addr_r[1]), .O(n16189));
    defparam rd_addr_r_0__bdd_4_lut_13795.LUT_INIT = 16'he4aa;
    SB_LUT4 i4546_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_13_6 ), .O(n6020));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4546_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4545_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_13_5 ), .O(n6019));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4545_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16189_bdd_4_lut (.I0(n16189), .I1(\REG.mem_21_31 ), .I2(\REG.mem_20_31 ), 
            .I3(rd_addr_r[1]), .O(n16192));
    defparam n16189_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12543 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_23 ), 
            .I2(\REG.mem_7_23 ), .I3(rd_addr_r[1]), .O(n14665));
    defparam rd_addr_r_0__bdd_4_lut_12543.LUT_INIT = 16'he4aa;
    SB_LUT4 n14665_bdd_4_lut (.I0(n14665), .I1(\REG.mem_5_23 ), .I2(\REG.mem_4_23 ), 
            .I3(rd_addr_r[1]), .O(n14668));
    defparam n14665_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12587 (.I0(rd_addr_r[1]), .I1(n13099), 
            .I2(n13100), .I3(rd_addr_r[2]), .O(n14659));
    defparam rd_addr_r_1__bdd_4_lut_12587.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13131 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_6 ), 
            .I2(\REG.mem_11_6 ), .I3(rd_addr_r[1]), .O(n15391));
    defparam rd_addr_r_0__bdd_4_lut_13131.LUT_INIT = 16'he4aa;
    SB_DFF i1151_1152 (.Q(\REG.mem_11_19 ), .C(FIFO_CLK_c), .D(n5969));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n15391_bdd_4_lut (.I0(n15391), .I1(\REG.mem_9_6 ), .I2(\REG.mem_8_6 ), 
            .I3(rd_addr_r[1]), .O(n13929));
    defparam n15391_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR wr_grey_sync_r__i2 (.Q(\wr_grey_sync_r[2] ), .C(FIFO_CLK_c), 
            .D(wr_grey_w[2]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_LUT4 n14659_bdd_4_lut (.I0(n14659), .I1(n13091), .I2(n13090), .I3(rd_addr_r[2]), 
            .O(n14662));
    defparam n14659_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut (.I0(rd_addr_r[1]), .I1(n14116), .I2(n14117), 
            .I3(rd_addr_r[2]), .O(n16183));
    defparam rd_addr_r_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n16183_bdd_4_lut (.I0(n16183), .I1(n14111), .I2(n14110), .I3(rd_addr_r[2]), 
            .O(n13568));
    defparam n16183_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR wr_grey_sync_r__i3 (.Q(\wr_grey_sync_r[3] ), .C(FIFO_CLK_c), 
            .D(wr_grey_w[3]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFSR wr_grey_sync_r__i4 (.Q(\wr_grey_sync_r[4] ), .C(FIFO_CLK_c), 
            .D(wr_grey_w[4]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFF i1148_1149 (.Q(\REG.mem_11_18 ), .C(FIFO_CLK_c), .D(n5968));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1145_1146 (.Q(\REG.mem_11_17 ), .C(FIFO_CLK_c), .D(n5967));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1142_1143 (.Q(\REG.mem_11_16 ), .C(FIFO_CLK_c), .D(n5966));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1139_1140 (.Q(\REG.mem_11_15 ), .C(FIFO_CLK_c), .D(n5965));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1136_1137 (.Q(\REG.mem_11_14 ), .C(FIFO_CLK_c), .D(n5964));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12528 (.I0(rd_addr_r[2]), .I1(n13167), 
            .I2(n13170), .I3(rd_addr_r[3]), .O(n14653));
    defparam rd_addr_r_2__bdd_4_lut_12528.LUT_INIT = 16'he4aa;
    SB_LUT4 i4138_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_0_31 ), .O(n5612));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4138_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13790 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_30 ), 
            .I2(\REG.mem_15_30 ), .I3(rd_addr_r[1]), .O(n16177));
    defparam rd_addr_r_0__bdd_4_lut_13790.LUT_INIT = 16'he4aa;
    SB_LUT4 n16177_bdd_4_lut (.I0(n16177), .I1(\REG.mem_13_30 ), .I2(\REG.mem_12_30 ), 
            .I3(rd_addr_r[1]), .O(n16180));
    defparam n16177_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14653_bdd_4_lut (.I0(n14653), .I1(n13164), .I2(n13161), .I3(rd_addr_r[3]), 
            .O(n14656));
    defparam n14653_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12518 (.I0(rd_addr_r[1]), .I1(n13069), 
            .I2(n13070), .I3(rd_addr_r[2]), .O(n14647));
    defparam rd_addr_r_1__bdd_4_lut_12518.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13181 (.I0(rd_addr_r[1]), .I1(n13411), 
            .I2(n13412), .I3(rd_addr_r[2]), .O(n15385));
    defparam rd_addr_r_1__bdd_4_lut_13181.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_r_5__I_0_123_i1_3_lut (.I0(\wr_addr_r[0] ), .I1(\wr_addr_p1_w[0] ), 
            .I2(wr_fifo_en_w), .I3(GND_net), .O(wr_addr_nxt_c[0]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_5__I_0_123_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13780 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_31 ), 
            .I2(\REG.mem_27_31 ), .I3(rd_addr_r[1]), .O(n16171));
    defparam rd_addr_r_0__bdd_4_lut_13780.LUT_INIT = 16'he4aa;
    SB_DFF i1133_1134 (.Q(\REG.mem_11_13 ), .C(FIFO_CLK_c), .D(n5963));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1130_1131 (.Q(\REG.mem_11_12 ), .C(FIFO_CLK_c), .D(n5962));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n16171_bdd_4_lut (.I0(n16171), .I1(\REG.mem_25_31 ), .I2(\REG.mem_24_31 ), 
            .I3(rd_addr_r[1]), .O(n16174));
    defparam n16171_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15385_bdd_4_lut (.I0(n15385), .I1(n13406), .I2(n13405), .I3(rd_addr_r[2]), 
            .O(n13445));
    defparam n15385_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1127_1128 (.Q(\REG.mem_11_11 ), .C(FIFO_CLK_c), .D(n5961));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1124_1125 (.Q(\REG.mem_11_10 ), .C(FIFO_CLK_c), .D(n5960));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1121_1122 (.Q(\REG.mem_11_9 ), .C(FIFO_CLK_c), .D(n5959));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1118_1119 (.Q(\REG.mem_11_8 ), .C(FIFO_CLK_c), .D(n5958));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1115_1116 (.Q(\REG.mem_11_7 ), .C(FIFO_CLK_c), .D(n5957));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1112_1113 (.Q(\REG.mem_11_6 ), .C(FIFO_CLK_c), .D(n5956));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1109_1110 (.Q(\REG.mem_11_5 ), .C(FIFO_CLK_c), .D(n5955));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1106_1107 (.Q(\REG.mem_11_4 ), .C(FIFO_CLK_c), .D(n5954));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1103_1104 (.Q(\REG.mem_11_3 ), .C(FIFO_CLK_c), .D(n5953));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_13261 (.I0(rd_addr_r[3]), .I1(n13609), 
            .I2(n13610), .I3(rd_addr_r[4]), .O(n15379));
    defparam rd_addr_r_3__bdd_4_lut_13261.LUT_INIT = 16'he4aa;
    SB_LUT4 n15379_bdd_4_lut (.I0(n15379), .I1(n13604), .I2(n15346), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[12]));
    defparam n15379_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4544_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_13_4 ), .O(n6018));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4544_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4543_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_13_3 ), .O(n6017));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4543_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_69 (.I0(wp_sync2_r[5]), .I1(wp_sync2_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n4814));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_69.LUT_INIT = 16'h6666;
    SB_LUT4 i4139_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_0_30 ), .O(n5613));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4139_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_13815 (.I0(rd_addr_r[2]), .I1(n15052), 
            .I2(n14602), .I3(rd_addr_r[3]), .O(n16153));
    defparam rd_addr_r_2__bdd_4_lut_13815.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12428 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_22 ), 
            .I2(\REG.mem_11_22 ), .I3(rd_addr_r[1]), .O(n14545));
    defparam rd_addr_r_0__bdd_4_lut_12428.LUT_INIT = 16'he4aa;
    SB_LUT4 n16153_bdd_4_lut (.I0(n16153), .I1(n15226), .I2(n15322), .I3(rd_addr_r[3]), 
            .O(n16156));
    defparam n16153_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13775 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_31 ), 
            .I2(\REG.mem_31_31 ), .I3(rd_addr_r[1]), .O(n16147));
    defparam rd_addr_r_0__bdd_4_lut_13775.LUT_INIT = 16'he4aa;
    SB_DFF i1100_1101 (.Q(\REG.mem_11_2 ), .C(FIFO_CLK_c), .D(n5952));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1097_1098 (.Q(\REG.mem_11_1 ), .C(FIFO_CLK_c), .D(n5951));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1094_1095 (.Q(\REG.mem_11_0 ), .C(FIFO_CLK_c), .D(n5950));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1091_1092 (.Q(\REG.mem_10_31 ), .C(FIFO_CLK_c), .D(n5949));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1088_1089 (.Q(\REG.mem_10_30 ), .C(FIFO_CLK_c), .D(n5948));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1085_1086 (.Q(\REG.mem_10_29 ), .C(FIFO_CLK_c), .D(n5947));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1082_1083 (.Q(\REG.mem_10_28 ), .C(FIFO_CLK_c), .D(n5946));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1079_1080 (.Q(\REG.mem_10_27 ), .C(FIFO_CLK_c), .D(n5945));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i128_129 (.Q(\REG.mem_0_30 ), .C(FIFO_CLK_c), .D(n5613));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13126 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_13 ), 
            .I2(\REG.mem_31_13 ), .I3(rd_addr_r[1]), .O(n15367));
    defparam rd_addr_r_0__bdd_4_lut_13126.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_70 (.I0(wp_sync2_r[0]), .I1(wp_sync_w[1]), .I2(GND_net), 
            .I3(GND_net), .O(wp_sync_w[0]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_70.LUT_INIT = 16'h6666;
    SB_LUT4 n15367_bdd_4_lut (.I0(n15367), .I1(\REG.mem_29_13 ), .I2(\REG.mem_28_13 ), 
            .I3(rd_addr_r[1]), .O(n13932));
    defparam n15367_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_71 (.I0(wp_sync2_r[2]), .I1(wp_sync_w[3]), .I2(GND_net), 
            .I3(GND_net), .O(wp_sync_w[2]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_71.LUT_INIT = 16'h6666;
    SB_LUT4 n14545_bdd_4_lut (.I0(n14545), .I1(\REG.mem_9_22 ), .I2(\REG.mem_8_22 ), 
            .I3(rd_addr_r[1]), .O(n14548));
    defparam n14545_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10853_4_lut (.I0(rd_addr_r[3]), .I1(rd_addr_r[0]), .I2(wp_sync_w[3]), 
            .I3(wp_sync_w[0]), .O(n12960));
    defparam i10853_4_lut.LUT_INIT = 16'h7bde;
    SB_DFF i131_132 (.Q(\REG.mem_0_31 ), .C(FIFO_CLK_c), .D(n5612));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1076_1077 (.Q(\REG.mem_10_26 ), .C(FIFO_CLK_c), .D(n5944));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i2_4_lut_adj_72 (.I0(wp_sync2_r[5]), .I1(rd_addr_p1_w[1]), .I2(rd_addr_p1_w[5]), 
            .I3(wp_sync_w[1]), .O(n8_adj_1387));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i2_4_lut_adj_72.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut (.I0(rd_addr_p1_w[2]), .I1(rd_addr_p1_w[0]), .I2(wp_sync_w[2]), 
            .I3(wp_sync_w[0]), .O(n7_adj_1388));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i1_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 n16147_bdd_4_lut (.I0(n16147), .I1(\REG.mem_29_31 ), .I2(\REG.mem_28_31 ), 
            .I3(rd_addr_r[1]), .O(n16150));
    defparam n16147_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4667_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_16_31 ), .O(n6141));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4667_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4666_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_16_30 ), .O(n6140));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4666_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14581_bdd_4_lut (.I0(n14581), .I1(\REG.mem_1_18 ), .I2(\REG.mem_0_18 ), 
            .I3(rd_addr_r[1]), .O(n14584));
    defparam n14581_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1073_1074 (.Q(\REG.mem_10_25 ), .C(FIFO_CLK_c), .D(n5943));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1070_1071 (.Q(\REG.mem_10_24 ), .C(FIFO_CLK_c), .D(n5942));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i215_216 (.Q(\REG.mem_1_27 ), .C(FIFO_CLK_c), .D(n5611));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3_4_lut (.I0(rd_addr_p1_w[3]), .I1(rd_addr_p1_w[4]), .I2(wp_sync_w[3]), 
            .I3(n4814), .O(n9_c));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i3_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13785 (.I0(rd_addr_r[1]), .I1(n13552), 
            .I2(n13553), .I3(rd_addr_r[2]), .O(n16141));
    defparam rd_addr_r_1__bdd_4_lut_13785.LUT_INIT = 16'he4aa;
    SB_LUT4 n16141_bdd_4_lut (.I0(n16141), .I1(n13544), .I2(n13543), .I3(rd_addr_r[2]), 
            .O(n13583));
    defparam n16141_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4665_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_16_29 ), .O(n6139));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4665_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13121 (.I0(rd_addr_r[1]), .I1(n13654), 
            .I2(n13655), .I3(rd_addr_r[2]), .O(n15361));
    defparam rd_addr_r_1__bdd_4_lut_13121.LUT_INIT = 16'he4aa;
    SB_LUT4 i4664_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_16_28 ), .O(n6138));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4664_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut (.I0(n12960), .I1(rd_addr_r[2]), .I2(dc32_fifo_empty), 
            .I3(wp_sync_w[2]), .O(n10_adj_1389));
    defparam i4_4_lut.LUT_INIT = 16'h4010;
    SB_LUT4 i5_3_lut (.I0(n9_c), .I1(n7_adj_1388), .I2(n8_adj_1387), .I3(GND_net), 
            .O(n12277));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4663_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_16_27 ), .O(n6137));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4663_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4662_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_16_26 ), .O(n6136));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4662_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4661_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_16_25 ), .O(n6135));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4661_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10907_4_lut (.I0(rd_addr_r[4]), .I1(rd_addr_r[1]), .I2(n4814), 
            .I3(wp_sync_w[1]), .O(n13016));
    defparam i10907_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 empty_nxt_c_I_11_4_lut (.I0(n13016), .I1(n12277), .I2(rd_fifo_en_w), 
            .I3(n10_adj_1389), .O(empty_nxt_c_N_636));   // src/fifo_dc_32_lut_gen.v(555[46:103])
    defparam empty_nxt_c_I_11_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 n15361_bdd_4_lut (.I0(n15361), .I1(n13799), .I2(n13798), .I3(rd_addr_r[2]), 
            .O(n15364));
    defparam n15361_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11004_3_lut (.I0(\REG.mem_22_17 ), .I1(\REG.mem_23_17 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13115));
    defparam i11004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13750 (.I0(rd_addr_r[1]), .I1(n14125), 
            .I2(n14126), .I3(rd_addr_r[2]), .O(n16135));
    defparam rd_addr_r_1__bdd_4_lut_13750.LUT_INIT = 16'he4aa;
    SB_LUT4 i4660_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_16_24 ), .O(n6134));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4660_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11003_3_lut (.I0(\REG.mem_20_17 ), .I1(\REG.mem_21_17 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13114));
    defparam i11003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_5__I_0_i2_3_lut (.I0(rd_addr_r[1]), .I1(rd_addr_p1_w[1]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_5__N_573[1] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_5__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n16135_bdd_4_lut (.I0(n16135), .I1(n14120), .I2(n14119), .I3(rd_addr_r[2]), 
            .O(n14159));
    defparam n16135_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4659_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_16_23 ), .O(n6133));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4659_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13755 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_15 ), 
            .I2(\REG.mem_23_15 ), .I3(rd_addr_r[1]), .O(n16129));
    defparam rd_addr_r_0__bdd_4_lut_13755.LUT_INIT = 16'he4aa;
    SB_LUT4 i4658_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_16_22 ), .O(n6132));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4658_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4657_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_16_21 ), .O(n6131));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4657_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4656_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_16_20 ), .O(n6130));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4656_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4542_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_13_2 ), .O(n6016));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4542_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16129_bdd_4_lut (.I0(n16129), .I1(\REG.mem_21_15 ), .I2(\REG.mem_20_15 ), 
            .I3(rd_addr_r[1]), .O(n16132));
    defparam n16129_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4655_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_16_19 ), .O(n6129));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4655_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13106 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_24 ), 
            .I2(\REG.mem_7_24 ), .I3(rd_addr_r[1]), .O(n15355));
    defparam rd_addr_r_0__bdd_4_lut_13106.LUT_INIT = 16'he4aa;
    SB_LUT4 i4654_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_16_18 ), .O(n6128));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4654_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4653_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_16_17 ), .O(n6127));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4653_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15355_bdd_4_lut (.I0(n15355), .I1(\REG.mem_5_24 ), .I2(\REG.mem_4_24 ), 
            .I3(rd_addr_r[1]), .O(n13935));
    defparam n15355_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13096 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_6 ), 
            .I2(\REG.mem_15_6 ), .I3(rd_addr_r[1]), .O(n15349));
    defparam rd_addr_r_0__bdd_4_lut_13096.LUT_INIT = 16'he4aa;
    SB_LUT4 i4652_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_16_16 ), .O(n6126));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4652_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15349_bdd_4_lut (.I0(n15349), .I1(\REG.mem_13_6 ), .I2(\REG.mem_12_6 ), 
            .I3(rd_addr_r[1]), .O(n13938));
    defparam n15349_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4651_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_16_15 ), .O(n6125));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4651_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4650_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_16_14 ), .O(n6124));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4650_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13740 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_4 ), 
            .I2(\REG.mem_3_4 ), .I3(rd_addr_r[1]), .O(n16111));
    defparam rd_addr_r_0__bdd_4_lut_13740.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13101 (.I0(rd_addr_r[1]), .I1(n13717), 
            .I2(n13718), .I3(rd_addr_r[2]), .O(n15343));
    defparam rd_addr_r_1__bdd_4_lut_13101.LUT_INIT = 16'he4aa;
    SB_LUT4 n15343_bdd_4_lut (.I0(n15343), .I1(n13439), .I2(n13438), .I3(rd_addr_r[2]), 
            .O(n15346));
    defparam n15343_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16111_bdd_4_lut (.I0(n16111), .I1(\REG.mem_1_4 ), .I2(\REG.mem_0_4 ), 
            .I3(rd_addr_r[1]), .O(n16114));
    defparam n16111_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4541_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_13_1 ), .O(n6015));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4541_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4649_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_16_13 ), .O(n6123));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4649_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4540_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_13_0 ), .O(n6014));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4540_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4648_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_16_12 ), .O(n6122));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4648_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4647_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_16_11 ), .O(n6121));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4647_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4646_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_16_10 ), .O(n6120));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4646_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4645_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_16_9 ), .O(n6119));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4645_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4644_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_16_8 ), .O(n6118));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4644_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4643_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_16_7 ), .O(n6117));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4643_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13745 (.I0(rd_addr_r[1]), .I1(n13195), 
            .I2(n13196), .I3(rd_addr_r[2]), .O(n16105));
    defparam rd_addr_r_1__bdd_4_lut_13745.LUT_INIT = 16'he4aa;
    SB_LUT4 i4642_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_16_6 ), .O(n6116));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4642_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4641_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_16_5 ), .O(n6115));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4641_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4640_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_16_4 ), .O(n6114));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4640_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16105_bdd_4_lut (.I0(n16105), .I1(n13193), .I2(n13192), .I3(rd_addr_r[2]), 
            .O(n13211));
    defparam n16105_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4639_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_16_3 ), .O(n6113));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4639_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_13236 (.I0(rd_addr_r[2]), .I1(n13887), 
            .I2(n13902), .I3(rd_addr_r[3]), .O(n15337));
    defparam rd_addr_r_2__bdd_4_lut_13236.LUT_INIT = 16'he4aa;
    SB_LUT4 i4140_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_0_29 ), .O(n5614));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4140_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_13760 (.I0(rd_addr_r[2]), .I1(n14770), 
            .I2(n14758), .I3(rd_addr_r[3]), .O(n16099));
    defparam rd_addr_r_2__bdd_4_lut_13760.LUT_INIT = 16'he4aa;
    SB_LUT4 n15337_bdd_4_lut (.I0(n15337), .I1(n13884), .I2(n13869), .I3(rd_addr_r[3]), 
            .O(n15340));
    defparam n15337_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5051_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_28_31 ), .O(n6525));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5051_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16099_bdd_4_lut (.I0(n16099), .I1(n14914), .I2(n14926), .I3(rd_addr_r[3]), 
            .O(n16102));
    defparam n16099_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13091 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_24 ), 
            .I2(\REG.mem_11_24 ), .I3(rd_addr_r[1]), .O(n15331));
    defparam rd_addr_r_0__bdd_4_lut_13091.LUT_INIT = 16'he4aa;
    SB_LUT4 i4638_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_16_2 ), .O(n6112));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4638_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4637_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_16_1 ), .O(n6111));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4637_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15331_bdd_4_lut (.I0(n15331), .I1(\REG.mem_9_24 ), .I2(\REG.mem_8_24 ), 
            .I3(rd_addr_r[1]), .O(n13944));
    defparam n15331_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4636_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_16_0 ), .O(n6110));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4636_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13720 (.I0(rd_addr_r[1]), .I1(n13576), 
            .I2(n13577), .I3(rd_addr_r[2]), .O(n16087));
    defparam rd_addr_r_1__bdd_4_lut_13720.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13076 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_28 ), 
            .I2(\REG.mem_23_28 ), .I3(rd_addr_r[1]), .O(n15325));
    defparam rd_addr_r_0__bdd_4_lut_13076.LUT_INIT = 16'he4aa;
    SB_LUT4 n15325_bdd_4_lut (.I0(n15325), .I1(\REG.mem_21_28 ), .I2(\REG.mem_20_28 ), 
            .I3(rd_addr_r[1]), .O(n13947));
    defparam n15325_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16087_bdd_4_lut (.I0(n16087), .I1(n13550), .I2(n13549), .I3(rd_addr_r[2]), 
            .O(n13610));
    defparam n16087_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13071 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_21 ), 
            .I2(\REG.mem_19_21 ), .I3(rd_addr_r[1]), .O(n15319));
    defparam rd_addr_r_0__bdd_4_lut_13071.LUT_INIT = 16'he4aa;
    SB_LUT4 n15319_bdd_4_lut (.I0(n15319), .I1(\REG.mem_17_21 ), .I2(\REG.mem_16_21 ), 
            .I3(rd_addr_r[1]), .O(n15322));
    defparam n15319_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5050_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_28_30 ), .O(n6524));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5050_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13725 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_24 ), 
            .I2(\REG.mem_31_24 ), .I3(rd_addr_r[1]), .O(n16075));
    defparam rd_addr_r_0__bdd_4_lut_13725.LUT_INIT = 16'he4aa;
    SB_LUT4 n16075_bdd_4_lut (.I0(n16075), .I1(\REG.mem_29_24 ), .I2(\REG.mem_28_24 ), 
            .I3(rd_addr_r[1]), .O(n13614));
    defparam n16075_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13066 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_0 ), 
            .I2(\REG.mem_7_0 ), .I3(rd_addr_r[1]), .O(n15313));
    defparam rd_addr_r_0__bdd_4_lut_13066.LUT_INIT = 16'he4aa;
    SB_LUT4 n15313_bdd_4_lut (.I0(n15313), .I1(\REG.mem_5_0 ), .I2(\REG.mem_4_0 ), 
            .I3(rd_addr_r[1]), .O(n13452));
    defparam n15313_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12453 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_4 ), 
            .I2(\REG.mem_11_4 ), .I3(rd_addr_r[1]), .O(n14575));
    defparam rd_addr_r_0__bdd_4_lut_12453.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13086 (.I0(rd_addr_r[1]), .I1(n13135), 
            .I2(n13136), .I3(rd_addr_r[2]), .O(n15307));
    defparam rd_addr_r_1__bdd_4_lut_13086.LUT_INIT = 16'he4aa;
    SB_DFF i188_189 (.Q(\REG.mem_1_18 ), .C(FIFO_CLK_c), .D(n5610));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1067_1068 (.Q(\REG.mem_10_23 ), .C(FIFO_CLK_c), .D(n5941));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1064_1065 (.Q(\REG.mem_10_22 ), .C(FIFO_CLK_c), .D(n5940));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1061_1062 (.Q(\REG.mem_10_21 ), .C(FIFO_CLK_c), .D(n5939));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1058_1059 (.Q(\REG.mem_10_20 ), .C(FIFO_CLK_c), .D(n5938));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1055_1056 (.Q(\REG.mem_10_19 ), .C(FIFO_CLK_c), .D(n5937));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i203_204 (.Q(\REG.mem_1_23 ), .C(FIFO_CLK_c), .D(n5608));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i134_135 (.Q(\REG.mem_1_0 ), .C(FIFO_CLK_c), .D(n5604));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5049_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_28_29 ), .O(n6523));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5049_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15307_bdd_4_lut (.I0(n15307), .I1(n13127), .I2(n13126), .I3(rd_addr_r[2]), 
            .O(n13454));
    defparam n15307_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_13081 (.I0(rd_addr_r[2]), .I1(n13917), 
            .I2(n13932), .I3(rd_addr_r[3]), .O(n15301));
    defparam rd_addr_r_2__bdd_4_lut_13081.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13695 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_27 ), 
            .I2(\REG.mem_27_27 ), .I3(rd_addr_r[1]), .O(n16057));
    defparam rd_addr_r_0__bdd_4_lut_13695.LUT_INIT = 16'he4aa;
    SB_LUT4 n16057_bdd_4_lut (.I0(n16057), .I1(\REG.mem_25_27 ), .I2(\REG.mem_24_27 ), 
            .I3(rd_addr_r[1]), .O(n16060));
    defparam n16057_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15301_bdd_4_lut (.I0(n15301), .I1(n13914), .I2(n13641), .I3(rd_addr_r[3]), 
            .O(n15304));
    defparam n15301_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i137_138 (.Q(\REG.mem_1_1 ), .C(FIFO_CLK_c), .D(n5603));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i140_141 (.Q(\REG.mem_1_2 ), .C(FIFO_CLK_c), .D(n5602));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i38_39 (.Q(\REG.mem_0_0 ), .C(FIFO_CLK_c), .D(n5601));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1052_1053 (.Q(\REG.mem_10_18 ), .C(FIFO_CLK_c), .D(n5936));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13061 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_6 ), 
            .I2(\REG.mem_19_6 ), .I3(rd_addr_r[1]), .O(n15295));
    defparam rd_addr_r_0__bdd_4_lut_13061.LUT_INIT = 16'he4aa;
    SB_LUT4 i5048_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_28_28 ), .O(n6522));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5048_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5047_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_28_27 ), .O(n6521));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5047_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13680 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_24 ), 
            .I2(\REG.mem_19_24 ), .I3(rd_addr_r[1]), .O(n16051));
    defparam rd_addr_r_0__bdd_4_lut_13680.LUT_INIT = 16'he4aa;
    SB_LUT4 i5046_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_28_26 ), .O(n6520));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5046_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15295_bdd_4_lut (.I0(n15295), .I1(\REG.mem_17_6 ), .I2(\REG.mem_16_6 ), 
            .I3(rd_addr_r[1]), .O(n13953));
    defparam n15295_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16051_bdd_4_lut (.I0(n16051), .I1(\REG.mem_17_24 ), .I2(\REG.mem_16_24 ), 
            .I3(rd_addr_r[1]), .O(n13629));
    defparam n16051_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1049_1050 (.Q(\REG.mem_10_17 ), .C(FIFO_CLK_c), .D(n5935));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1046_1047 (.Q(\REG.mem_10_16 ), .C(FIFO_CLK_c), .D(n5934));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1043_1044 (.Q(\REG.mem_10_15 ), .C(FIFO_CLK_c), .D(n5933));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4142_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_0_28 ), .O(n5616));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4142_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5045_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_28_25 ), .O(n6519));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5045_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5044_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_28_24 ), .O(n6518));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5044_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5043_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_28_23 ), .O(n6517));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5043_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13046 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_24 ), 
            .I2(\REG.mem_15_24 ), .I3(rd_addr_r[1]), .O(n15289));
    defparam rd_addr_r_0__bdd_4_lut_13046.LUT_INIT = 16'he4aa;
    SB_LUT4 i11180_3_lut (.I0(\REG.mem_0_17 ), .I1(\REG.mem_1_17 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13291));
    defparam i11180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11181_3_lut (.I0(\REG.mem_2_17 ), .I1(\REG.mem_3_17 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13292));
    defparam i11181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n14575_bdd_4_lut (.I0(n14575), .I1(\REG.mem_9_4 ), .I2(\REG.mem_8_4 ), 
            .I3(rd_addr_r[1]), .O(n14578));
    defparam n14575_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4143_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_0_27 ), .O(n5617));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4143_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15289_bdd_4_lut (.I0(n15289), .I1(\REG.mem_13_24 ), .I2(\REG.mem_12_24 ), 
            .I3(rd_addr_r[1]), .O(n13956));
    defparam n15289_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4146_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_0_26 ), .O(n5620));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4146_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5042_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_28_22 ), .O(n6516));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5042_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4147_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_0_25 ), .O(n5621));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4147_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13675 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_8 ), 
            .I2(\REG.mem_23_8 ), .I3(rd_addr_r[1]), .O(n16039));
    defparam rd_addr_r_0__bdd_4_lut_13675.LUT_INIT = 16'he4aa;
    SB_LUT4 i5041_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_28_21 ), .O(n6515));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5041_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5040_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_28_20 ), .O(n6514));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5040_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11199_3_lut (.I0(\REG.mem_6_17 ), .I1(\REG.mem_7_17 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13310));
    defparam i11199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11198_3_lut (.I0(\REG.mem_4_17 ), .I1(\REG.mem_5_17 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13309));
    defparam i11198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n16039_bdd_4_lut (.I0(n16039), .I1(\REG.mem_21_8 ), .I2(\REG.mem_20_8 ), 
            .I3(rd_addr_r[1]), .O(n13632));
    defparam n16039_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5039_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_28_19 ), .O(n6513));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5039_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_13116 (.I0(rd_addr_r[3]), .I1(n13054), 
            .I2(n13055), .I3(rd_addr_r[4]), .O(n15277));
    defparam rd_addr_r_3__bdd_4_lut_13116.LUT_INIT = 16'he4aa;
    SB_LUT4 n15277_bdd_4_lut (.I0(n15277), .I1(n13583), .I2(n13582), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[31]));
    defparam n15277_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_73 (.I0(dc32_fifo_empty), .I1(dc32_fifo_read_enable), 
            .I2(GND_net), .I3(GND_net), .O(rd_fifo_en_w));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i1_2_lut_adj_73.LUT_INIT = 16'h4444;
    SB_LUT4 i10992_3_lut (.I0(n14788), .I1(n14752), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13103));
    defparam i10992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10993_3_lut (.I0(n14626), .I1(n13103), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n13104));
    defparam i10993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13041 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_16 ), 
            .I2(\REG.mem_23_16 ), .I3(rd_addr_r[1]), .O(n15271));
    defparam rd_addr_r_0__bdd_4_lut_13041.LUT_INIT = 16'he4aa;
    SB_LUT4 n15271_bdd_4_lut (.I0(n15271), .I1(\REG.mem_21_16 ), .I2(\REG.mem_20_16 ), 
            .I3(rd_addr_r[1]), .O(n15274));
    defparam n15271_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8141316_i1_3_lut (.I0(n14674), .I1(n13104), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[0]));
    defparam i8141316_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11249_3_lut (.I0(\REG.mem_16_2 ), .I1(\REG.mem_17_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13360));
    defparam i11249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13056 (.I0(rd_addr_r[1]), .I1(n13207), 
            .I2(n13208), .I3(rd_addr_r[2]), .O(n15265));
    defparam rd_addr_r_1__bdd_4_lut_13056.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_13715 (.I0(rd_addr_r[2]), .I1(n15586), 
            .I2(n15544), .I3(rd_addr_r[3]), .O(n16027));
    defparam rd_addr_r_2__bdd_4_lut_13715.LUT_INIT = 16'he4aa;
    SB_LUT4 i11250_3_lut (.I0(\REG.mem_18_2 ), .I1(\REG.mem_19_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13361));
    defparam i11250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n15265_bdd_4_lut (.I0(n15265), .I1(n13205), .I2(n13204), .I3(rd_addr_r[2]), 
            .O(n13964));
    defparam n15265_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5038_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_28_18 ), .O(n6512));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5038_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16027_bdd_4_lut (.I0(n16027), .I1(n15616), .I2(n15652), .I3(rd_addr_r[3]), 
            .O(n16030));
    defparam n16027_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5037_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_28_17 ), .O(n6511));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5037_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13026 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_6 ), 
            .I2(\REG.mem_23_6 ), .I3(rd_addr_r[1]), .O(n15253));
    defparam rd_addr_r_0__bdd_4_lut_13026.LUT_INIT = 16'he4aa;
    SB_LUT4 i11256_3_lut (.I0(\REG.mem_22_2 ), .I1(\REG.mem_23_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13367));
    defparam i11256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n15253_bdd_4_lut (.I0(n15253), .I1(\REG.mem_21_6 ), .I2(\REG.mem_20_6 ), 
            .I3(rd_addr_r[1]), .O(n13971));
    defparam n15253_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11255_3_lut (.I0(\REG.mem_20_2 ), .I1(\REG.mem_21_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13366));
    defparam i11255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13705 (.I0(rd_addr_r[1]), .I1(n13222), 
            .I2(n13223), .I3(rd_addr_r[2]), .O(n16021));
    defparam rd_addr_r_1__bdd_4_lut_13705.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13011 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_8 ), 
            .I2(\REG.mem_27_8 ), .I3(rd_addr_r[1]), .O(n15247));
    defparam rd_addr_r_0__bdd_4_lut_13011.LUT_INIT = 16'he4aa;
    SB_LUT4 n15247_bdd_4_lut (.I0(n15247), .I1(\REG.mem_25_8 ), .I2(\REG.mem_24_8 ), 
            .I3(rd_addr_r[1]), .O(n13974));
    defparam n15247_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5036_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_28_16 ), .O(n6510));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5036_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1040_1041 (.Q(\REG.mem_10_14 ), .C(FIFO_CLK_c), .D(n5932));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1037_1038 (.Q(\REG.mem_10_13 ), .C(FIFO_CLK_c), .D(n5931));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1034_1035 (.Q(\REG.mem_10_12 ), .C(FIFO_CLK_c), .D(n5930));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1031_1032 (.Q(\REG.mem_10_11 ), .C(FIFO_CLK_c), .D(n5929));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1028_1029 (.Q(\REG.mem_10_10 ), .C(FIFO_CLK_c), .D(n5928));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1025_1026 (.Q(\REG.mem_10_9 ), .C(FIFO_CLK_c), .D(n5927));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1022_1023 (.Q(\REG.mem_10_8 ), .C(FIFO_CLK_c), .D(n5926));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1019_1020 (.Q(\REG.mem_10_7 ), .C(FIFO_CLK_c), .D(n5925));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1016_1017 (.Q(\REG.mem_10_6 ), .C(FIFO_CLK_c), .D(n5924));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1013_1014 (.Q(\REG.mem_10_5 ), .C(FIFO_CLK_c), .D(n5923));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1010_1011 (.Q(\REG.mem_10_4 ), .C(FIFO_CLK_c), .D(n5922));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1007_1008 (.Q(\REG.mem_10_3 ), .C(FIFO_CLK_c), .D(n5921));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1004_1005 (.Q(\REG.mem_10_2 ), .C(FIFO_CLK_c), .D(n5920));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1001_1002 (.Q(\REG.mem_10_1 ), .C(FIFO_CLK_c), .D(n5919));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i998_999 (.Q(\REG.mem_10_0 ), .C(FIFO_CLK_c), .D(n5918));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i995_996 (.Q(\REG.mem_9_31 ), .C(FIFO_CLK_c), .D(n5917));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i992_993 (.Q(\REG.mem_9_30 ), .C(FIFO_CLK_c), .D(n5916));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i989_990 (.Q(\REG.mem_9_29 ), .C(FIFO_CLK_c), .D(n5915));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i986_987 (.Q(\REG.mem_9_28 ), .C(FIFO_CLK_c), .D(n5914));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i983_984 (.Q(\REG.mem_9_27 ), .C(FIFO_CLK_c), .D(n5913));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i980_981 (.Q(\REG.mem_9_26 ), .C(FIFO_CLK_c), .D(n5912));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i977_978 (.Q(\REG.mem_9_25 ), .C(FIFO_CLK_c), .D(n5911));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i974_975 (.Q(\REG.mem_9_24 ), .C(FIFO_CLK_c), .D(n5910));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i971_972 (.Q(\REG.mem_9_23 ), .C(FIFO_CLK_c), .D(n5909));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i968_969 (.Q(\REG.mem_9_22 ), .C(FIFO_CLK_c), .D(n5908));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i965_966 (.Q(\REG.mem_9_21 ), .C(FIFO_CLK_c), .D(n5907));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i962_963 (.Q(\REG.mem_9_20 ), .C(FIFO_CLK_c), .D(n5906));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i959_960 (.Q(\REG.mem_9_19 ), .C(FIFO_CLK_c), .D(n5905));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i956_957 (.Q(\REG.mem_9_18 ), .C(FIFO_CLK_c), .D(n5904));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i953_954 (.Q(\REG.mem_9_17 ), .C(FIFO_CLK_c), .D(n5903));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i950_951 (.Q(\REG.mem_9_16 ), .C(FIFO_CLK_c), .D(n5902));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i947_948 (.Q(\REG.mem_9_15 ), .C(FIFO_CLK_c), .D(n5901));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i944_945 (.Q(\REG.mem_9_14 ), .C(FIFO_CLK_c), .D(n5900));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i941_942 (.Q(\REG.mem_9_13 ), .C(FIFO_CLK_c), .D(n5899));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i938_939 (.Q(\REG.mem_9_12 ), .C(FIFO_CLK_c), .D(n5898));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i935_936 (.Q(\REG.mem_9_11 ), .C(FIFO_CLK_c), .D(n5897));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i932_933 (.Q(\REG.mem_9_10 ), .C(FIFO_CLK_c), .D(n5896));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i929_930 (.Q(\REG.mem_9_9 ), .C(FIFO_CLK_c), .D(n5895));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i926_927 (.Q(\REG.mem_9_8 ), .C(FIFO_CLK_c), .D(n5894));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i923_924 (.Q(\REG.mem_9_7 ), .C(FIFO_CLK_c), .D(n5893));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i920_921 (.Q(\REG.mem_9_6 ), .C(FIFO_CLK_c), .D(n5892));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i917_918 (.Q(\REG.mem_9_5 ), .C(FIFO_CLK_c), .D(n5891));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i914_915 (.Q(\REG.mem_9_4 ), .C(FIFO_CLK_c), .D(n5890));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i911_912 (.Q(\REG.mem_9_3 ), .C(FIFO_CLK_c), .D(n5889));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i908_909 (.Q(\REG.mem_9_2 ), .C(FIFO_CLK_c), .D(n5888));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i905_906 (.Q(\REG.mem_9_1 ), .C(FIFO_CLK_c), .D(n5887));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i902_903 (.Q(\REG.mem_9_0 ), .C(FIFO_CLK_c), .D(n5886));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i899_900 (.Q(\REG.mem_8_31 ), .C(FIFO_CLK_c), .D(n5885));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i896_897 (.Q(\REG.mem_8_30 ), .C(FIFO_CLK_c), .D(n5884));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i893_894 (.Q(\REG.mem_8_29 ), .C(FIFO_CLK_c), .D(n5883));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i890_891 (.Q(\REG.mem_8_28 ), .C(FIFO_CLK_c), .D(n5882));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i887_888 (.Q(\REG.mem_8_27 ), .C(FIFO_CLK_c), .D(n5881));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i884_885 (.Q(\REG.mem_8_26 ), .C(FIFO_CLK_c), .D(n5880));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i881_882 (.Q(\REG.mem_8_25 ), .C(FIFO_CLK_c), .D(n5879));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i878_879 (.Q(\REG.mem_8_24 ), .C(FIFO_CLK_c), .D(n5878));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i875_876 (.Q(\REG.mem_8_23 ), .C(FIFO_CLK_c), .D(n5877));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i872_873 (.Q(\REG.mem_8_22 ), .C(FIFO_CLK_c), .D(n5876));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i869_870 (.Q(\REG.mem_8_21 ), .C(FIFO_CLK_c), .D(n5875));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i866_867 (.Q(\REG.mem_8_20 ), .C(FIFO_CLK_c), .D(n5874));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i863_864 (.Q(\REG.mem_8_19 ), .C(FIFO_CLK_c), .D(n5873));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i860_861 (.Q(\REG.mem_8_18 ), .C(FIFO_CLK_c), .D(n5872));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i857_858 (.Q(\REG.mem_8_17 ), .C(FIFO_CLK_c), .D(n5871));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i854_855 (.Q(\REG.mem_8_16 ), .C(FIFO_CLK_c), .D(n5870));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i851_852 (.Q(\REG.mem_8_15 ), .C(FIFO_CLK_c), .D(n5869));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i848_849 (.Q(\REG.mem_8_14 ), .C(FIFO_CLK_c), .D(n5868));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i845_846 (.Q(\REG.mem_8_13 ), .C(FIFO_CLK_c), .D(n5867));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i842_843 (.Q(\REG.mem_8_12 ), .C(FIFO_CLK_c), .D(n5866));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i839_840 (.Q(\REG.mem_8_11 ), .C(FIFO_CLK_c), .D(n5865));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i836_837 (.Q(\REG.mem_8_10 ), .C(FIFO_CLK_c), .D(n5864));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i833_834 (.Q(\REG.mem_8_9 ), .C(FIFO_CLK_c), .D(n5863));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i830_831 (.Q(\REG.mem_8_8 ), .C(FIFO_CLK_c), .D(n5862));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i827_828 (.Q(\REG.mem_8_7 ), .C(FIFO_CLK_c), .D(n5861));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i824_825 (.Q(\REG.mem_8_6 ), .C(FIFO_CLK_c), .D(n5860));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i821_822 (.Q(\REG.mem_8_5 ), .C(FIFO_CLK_c), .D(n5859));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i818_819 (.Q(\REG.mem_8_4 ), .C(FIFO_CLK_c), .D(n5858));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i815_816 (.Q(\REG.mem_8_3 ), .C(FIFO_CLK_c), .D(n5857));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i812_813 (.Q(\REG.mem_8_2 ), .C(FIFO_CLK_c), .D(n5856));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i809_810 (.Q(\REG.mem_8_1 ), .C(FIFO_CLK_c), .D(n5855));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i806_807 (.Q(\REG.mem_8_0 ), .C(FIFO_CLK_c), .D(n5854));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i803_804 (.Q(\REG.mem_7_31 ), .C(FIFO_CLK_c), .D(n5853));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i800_801 (.Q(\REG.mem_7_30 ), .C(FIFO_CLK_c), .D(n5852));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i797_798 (.Q(\REG.mem_7_29 ), .C(FIFO_CLK_c), .D(n5851));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i794_795 (.Q(\REG.mem_7_28 ), .C(FIFO_CLK_c), .D(n5850));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i791_792 (.Q(\REG.mem_7_27 ), .C(FIFO_CLK_c), .D(n5849));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i788_789 (.Q(\REG.mem_7_26 ), .C(FIFO_CLK_c), .D(n5848));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i785_786 (.Q(\REG.mem_7_25 ), .C(FIFO_CLK_c), .D(n5847));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i782_783 (.Q(\REG.mem_7_24 ), .C(FIFO_CLK_c), .D(n5846));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i779_780 (.Q(\REG.mem_7_23 ), .C(FIFO_CLK_c), .D(n5845));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i776_777 (.Q(\REG.mem_7_22 ), .C(FIFO_CLK_c), .D(n5844));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i773_774 (.Q(\REG.mem_7_21 ), .C(FIFO_CLK_c), .D(n5843));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i770_771 (.Q(\REG.mem_7_20 ), .C(FIFO_CLK_c), .D(n5842));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i767_768 (.Q(\REG.mem_7_19 ), .C(FIFO_CLK_c), .D(n5841));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i764_765 (.Q(\REG.mem_7_18 ), .C(FIFO_CLK_c), .D(n5840));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i761_762 (.Q(\REG.mem_7_17 ), .C(FIFO_CLK_c), .D(n5839));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i758_759 (.Q(\REG.mem_7_16 ), .C(FIFO_CLK_c), .D(n5838));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i755_756 (.Q(\REG.mem_7_15 ), .C(FIFO_CLK_c), .D(n5837));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i752_753 (.Q(\REG.mem_7_14 ), .C(FIFO_CLK_c), .D(n5836));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i749_750 (.Q(\REG.mem_7_13 ), .C(FIFO_CLK_c), .D(n5835));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i746_747 (.Q(\REG.mem_7_12 ), .C(FIFO_CLK_c), .D(n5834));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i743_744 (.Q(\REG.mem_7_11 ), .C(FIFO_CLK_c), .D(n5833));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i740_741 (.Q(\REG.mem_7_10 ), .C(FIFO_CLK_c), .D(n5832));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i737_738 (.Q(\REG.mem_7_9 ), .C(FIFO_CLK_c), .D(n5831));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i734_735 (.Q(\REG.mem_7_8 ), .C(FIFO_CLK_c), .D(n5830));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i731_732 (.Q(\REG.mem_7_7 ), .C(FIFO_CLK_c), .D(n5829));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i728_729 (.Q(\REG.mem_7_6 ), .C(FIFO_CLK_c), .D(n5828));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i725_726 (.Q(\REG.mem_7_5 ), .C(FIFO_CLK_c), .D(n5827));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i722_723 (.Q(\REG.mem_7_4 ), .C(FIFO_CLK_c), .D(n5826));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i719_720 (.Q(\REG.mem_7_3 ), .C(FIFO_CLK_c), .D(n5825));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i716_717 (.Q(\REG.mem_7_2 ), .C(FIFO_CLK_c), .D(n5824));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i713_714 (.Q(\REG.mem_7_1 ), .C(FIFO_CLK_c), .D(n5823));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i710_711 (.Q(\REG.mem_7_0 ), .C(FIFO_CLK_c), .D(n5822));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i707_708 (.Q(\REG.mem_6_31 ), .C(FIFO_CLK_c), .D(n5821));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i704_705 (.Q(\REG.mem_6_30 ), .C(FIFO_CLK_c), .D(n5820));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i701_702 (.Q(\REG.mem_6_29 ), .C(FIFO_CLK_c), .D(n5819));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i698_699 (.Q(\REG.mem_6_28 ), .C(FIFO_CLK_c), .D(n5818));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i695_696 (.Q(\REG.mem_6_27 ), .C(FIFO_CLK_c), .D(n5817));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i692_693 (.Q(\REG.mem_6_26 ), .C(FIFO_CLK_c), .D(n5816));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i689_690 (.Q(\REG.mem_6_25 ), .C(FIFO_CLK_c), .D(n5815));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i686_687 (.Q(\REG.mem_6_24 ), .C(FIFO_CLK_c), .D(n5814));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i683_684 (.Q(\REG.mem_6_23 ), .C(FIFO_CLK_c), .D(n5813));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i680_681 (.Q(\REG.mem_6_22 ), .C(FIFO_CLK_c), .D(n5812));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i677_678 (.Q(\REG.mem_6_21 ), .C(FIFO_CLK_c), .D(n5811));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i674_675 (.Q(\REG.mem_6_20 ), .C(FIFO_CLK_c), .D(n5810));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i671_672 (.Q(\REG.mem_6_19 ), .C(FIFO_CLK_c), .D(n5809));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i668_669 (.Q(\REG.mem_6_18 ), .C(FIFO_CLK_c), .D(n5808));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i665_666 (.Q(\REG.mem_6_17 ), .C(FIFO_CLK_c), .D(n5807));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i662_663 (.Q(\REG.mem_6_16 ), .C(FIFO_CLK_c), .D(n5806));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i659_660 (.Q(\REG.mem_6_15 ), .C(FIFO_CLK_c), .D(n5805));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i656_657 (.Q(\REG.mem_6_14 ), .C(FIFO_CLK_c), .D(n5804));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i653_654 (.Q(\REG.mem_6_13 ), .C(FIFO_CLK_c), .D(n5803));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i650_651 (.Q(\REG.mem_6_12 ), .C(FIFO_CLK_c), .D(n5802));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i647_648 (.Q(\REG.mem_6_11 ), .C(FIFO_CLK_c), .D(n5801));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i644_645 (.Q(\REG.mem_6_10 ), .C(FIFO_CLK_c), .D(n5800));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i641_642 (.Q(\REG.mem_6_9 ), .C(FIFO_CLK_c), .D(n5799));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i638_639 (.Q(\REG.mem_6_8 ), .C(FIFO_CLK_c), .D(n5798));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i635_636 (.Q(\REG.mem_6_7 ), .C(FIFO_CLK_c), .D(n5797));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i632_633 (.Q(\REG.mem_6_6 ), .C(FIFO_CLK_c), .D(n5796));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i629_630 (.Q(\REG.mem_6_5 ), .C(FIFO_CLK_c), .D(n5795));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i626_627 (.Q(\REG.mem_6_4 ), .C(FIFO_CLK_c), .D(n5794));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i623_624 (.Q(\REG.mem_6_3 ), .C(FIFO_CLK_c), .D(n5793));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i620_621 (.Q(\REG.mem_6_2 ), .C(FIFO_CLK_c), .D(n5792));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i617_618 (.Q(\REG.mem_6_1 ), .C(FIFO_CLK_c), .D(n5791));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i614_615 (.Q(\REG.mem_6_0 ), .C(FIFO_CLK_c), .D(n5790));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i611_612 (.Q(\REG.mem_5_31 ), .C(FIFO_CLK_c), .D(n5789));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i608_609 (.Q(\REG.mem_5_30 ), .C(FIFO_CLK_c), .D(n5788));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i143_144 (.Q(\REG.mem_1_3 ), .C(FIFO_CLK_c), .D(n5600));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5035_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_28_15 ), .O(n6509));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5035_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i605_606 (.Q(\REG.mem_5_29 ), .C(FIFO_CLK_c), .D(n5787));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13006 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_27 ), 
            .I2(\REG.mem_31_27 ), .I3(rd_addr_r[1]), .O(n15241));
    defparam rd_addr_r_0__bdd_4_lut_13006.LUT_INIT = 16'he4aa;
    SB_LUT4 n15241_bdd_4_lut (.I0(n15241), .I1(\REG.mem_29_27 ), .I2(\REG.mem_28_27 ), 
            .I3(rd_addr_r[1]), .O(n15244));
    defparam n15241_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i53_2_lut_3_lut (.I0(n13_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n25_adj_5));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i53_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i52_2_lut_3_lut (.I0(n13_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n9));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i52_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i602_603 (.Q(\REG.mem_5_28 ), .C(FIFO_CLK_c), .D(n5786));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5034_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_28_14 ), .O(n6508));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5034_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4149_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_0_23 ), .O(n5623));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4149_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i599_600 (.Q(\REG.mem_5_27 ), .C(FIFO_CLK_c), .D(n5785));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5147_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_31_31 ), .O(n6621));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5147_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5033_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_28_13 ), .O(n6507));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5033_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16021_bdd_4_lut (.I0(n16021), .I1(n13220), .I2(n13219), .I3(rd_addr_r[2]), 
            .O(n13247));
    defparam n16021_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5146_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_31_30 ), .O(n6620));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5146_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i596_597 (.Q(\REG.mem_5_26 ), .C(FIFO_CLK_c), .D(n5784));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5145_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_31_29 ), .O(n6619));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5145_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5144_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_31_28 ), .O(n6618));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5144_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5143_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_31_27 ), .O(n6617));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5143_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5142_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_31_26 ), .O(n6616));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5142_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i593_594 (.Q(\REG.mem_5_25 ), .C(FIFO_CLK_c), .D(n5783));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5032_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_28_12 ), .O(n6506));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5032_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i590_591 (.Q(\REG.mem_5_24 ), .C(FIFO_CLK_c), .D(n5782));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5031_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_28_11 ), .O(n6505));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5031_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4150_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_0_22 ), .O(n5624));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4150_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13001 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_12 ), 
            .I2(\REG.mem_11_12 ), .I3(rd_addr_r[1]), .O(n15235));
    defparam rd_addr_r_0__bdd_4_lut_13001.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13665 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_20 ), 
            .I2(\REG.mem_11_20 ), .I3(rd_addr_r[1]), .O(n16015));
    defparam rd_addr_r_0__bdd_4_lut_13665.LUT_INIT = 16'he4aa;
    SB_LUT4 i5030_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_28_10 ), .O(n6504));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5030_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_en_i_I_0_2_lut (.I0(dc32_fifo_write_enable), .I1(dc32_fifo_full), 
            .I2(GND_net), .I3(GND_net), .O(wr_fifo_en_w));   // src/fifo_dc_32_lut_gen.v(240[29:50])
    defparam wr_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 n16015_bdd_4_lut (.I0(n16015), .I1(\REG.mem_9_20 ), .I2(\REG.mem_8_20 ), 
            .I3(rd_addr_r[1]), .O(n16018));
    defparam n16015_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4151_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_0_21 ), .O(n5625));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4151_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5141_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_31_25 ), .O(n6615));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5141_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13646 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_13 ), 
            .I2(\REG.mem_19_13 ), .I3(rd_addr_r[1]), .O(n16009));
    defparam rd_addr_r_0__bdd_4_lut_13646.LUT_INIT = 16'he4aa;
    SB_LUT4 n16009_bdd_4_lut (.I0(n16009), .I1(\REG.mem_17_13 ), .I2(\REG.mem_16_13 ), 
            .I3(rd_addr_r[1]), .O(n13641));
    defparam n16009_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15235_bdd_4_lut (.I0(n15235), .I1(\REG.mem_9_12 ), .I2(\REG.mem_8_12 ), 
            .I3(rd_addr_r[1]), .O(n15238));
    defparam n15235_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5140_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_31_24 ), .O(n6614));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5140_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5139_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_31_23 ), .O(n6613));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5139_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5138_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_31_22 ), .O(n6612));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5138_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5029_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_28_9 ), .O(n6503));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5029_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5028_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_28_8 ), .O(n6502));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5028_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13641 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_16 ), 
            .I2(\REG.mem_3_16 ), .I3(rd_addr_r[1]), .O(n16003));
    defparam rd_addr_r_0__bdd_4_lut_13641.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12996 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_0 ), 
            .I2(\REG.mem_11_0 ), .I3(rd_addr_r[1]), .O(n15229));
    defparam rd_addr_r_0__bdd_4_lut_12996.LUT_INIT = 16'he4aa;
    SB_LUT4 n15229_bdd_4_lut (.I0(n15229), .I1(\REG.mem_9_0 ), .I2(\REG.mem_8_0 ), 
            .I3(rd_addr_r[1]), .O(n13464));
    defparam n15229_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5137_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_31_21 ), .O(n6611));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5137_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16003_bdd_4_lut (.I0(n16003), .I1(\REG.mem_1_16 ), .I2(\REG.mem_0_16 ), 
            .I3(rd_addr_r[1]), .O(n13650));
    defparam n16003_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12991 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_21 ), 
            .I2(\REG.mem_23_21 ), .I3(rd_addr_r[1]), .O(n15223));
    defparam rd_addr_r_0__bdd_4_lut_12991.LUT_INIT = 16'he4aa;
    SB_LUT4 i5136_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_31_20 ), .O(n6610));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5136_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4154_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_0_20 ), .O(n5628));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4154_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13636 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_20 ), 
            .I2(\REG.mem_15_20 ), .I3(rd_addr_r[1]), .O(n15997));
    defparam rd_addr_r_0__bdd_4_lut_13636.LUT_INIT = 16'he4aa;
    SB_DFF i587_588 (.Q(\REG.mem_5_23 ), .C(FIFO_CLK_c), .D(n5781));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4096_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_0_1 ), .O(n5570));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4096_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15997_bdd_4_lut (.I0(n15997), .I1(\REG.mem_13_20 ), .I2(\REG.mem_12_20 ), 
            .I3(rd_addr_r[1]), .O(n16000));
    defparam n15997_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15223_bdd_4_lut (.I0(n15223), .I1(\REG.mem_21_21 ), .I2(\REG.mem_20_21 ), 
            .I3(rd_addr_r[1]), .O(n15226));
    defparam n15223_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i584_585 (.Q(\REG.mem_5_22 ), .C(FIFO_CLK_c), .D(n5780));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5027_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_28_7 ), .O(n6501));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5027_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5135_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_31_19 ), .O(n6609));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5135_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5134_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_31_18 ), .O(n6608));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5134_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13631 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_20 ), 
            .I2(\REG.mem_19_20 ), .I3(rd_addr_r[1]), .O(n15991));
    defparam rd_addr_r_0__bdd_4_lut_13631.LUT_INIT = 16'he4aa;
    SB_LUT4 n15991_bdd_4_lut (.I0(n15991), .I1(\REG.mem_17_20 ), .I2(\REG.mem_16_20 ), 
            .I3(rd_addr_r[1]), .O(n14226));
    defparam n15991_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5133_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_31_17 ), .O(n6607));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5133_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5132_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_31_16 ), .O(n6606));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5132_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5131_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_31_15 ), .O(n6605));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5131_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12986 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_1 ), 
            .I2(\REG.mem_11_1 ), .I3(rd_addr_r[1]), .O(n15217));
    defparam rd_addr_r_0__bdd_4_lut_12986.LUT_INIT = 16'he4aa;
    SB_LUT4 i5130_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_31_14 ), .O(n6604));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5130_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i581_582 (.Q(\REG.mem_5_21 ), .C(FIFO_CLK_c), .D(n5779));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n15217_bdd_4_lut (.I0(n15217), .I1(\REG.mem_9_1 ), .I2(\REG.mem_8_1 ), 
            .I3(rd_addr_r[1]), .O(n15220));
    defparam n15217_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i578_579 (.Q(\REG.mem_5_20 ), .C(FIFO_CLK_c), .D(n5778));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13626 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_20 ), 
            .I2(\REG.mem_23_20 ), .I3(rd_addr_r[1]), .O(n15979));
    defparam rd_addr_r_0__bdd_4_lut_13626.LUT_INIT = 16'he4aa;
    SB_LUT4 n15979_bdd_4_lut (.I0(n15979), .I1(\REG.mem_21_20 ), .I2(\REG.mem_20_20 ), 
            .I3(rd_addr_r[1]), .O(n14229));
    defparam n15979_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13616 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_20 ), 
            .I2(\REG.mem_27_20 ), .I3(rd_addr_r[1]), .O(n15973));
    defparam rd_addr_r_0__bdd_4_lut_13616.LUT_INIT = 16'he4aa;
    SB_LUT4 n15973_bdd_4_lut (.I0(n15973), .I1(\REG.mem_25_20 ), .I2(\REG.mem_24_20 ), 
            .I3(rd_addr_r[1]), .O(n14232));
    defparam n15973_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13611 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_25 ), 
            .I2(\REG.mem_23_25 ), .I3(rd_addr_r[1]), .O(n15967));
    defparam rd_addr_r_0__bdd_4_lut_13611.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12981 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_28 ), 
            .I2(\REG.mem_27_28 ), .I3(rd_addr_r[1]), .O(n15205));
    defparam rd_addr_r_0__bdd_4_lut_12981.LUT_INIT = 16'he4aa;
    SB_LUT4 n15205_bdd_4_lut (.I0(n15205), .I1(\REG.mem_25_28 ), .I2(\REG.mem_24_28 ), 
            .I3(rd_addr_r[1]), .O(n13980));
    defparam n15205_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i575_576 (.Q(\REG.mem_5_19 ), .C(FIFO_CLK_c), .D(n5777));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12971 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_30 ), 
            .I2(\REG.mem_11_30 ), .I3(rd_addr_r[1]), .O(n15199));
    defparam rd_addr_r_0__bdd_4_lut_12971.LUT_INIT = 16'he4aa;
    SB_LUT4 n15199_bdd_4_lut (.I0(n15199), .I1(\REG.mem_9_30 ), .I2(\REG.mem_8_30 ), 
            .I3(rd_addr_r[1]), .O(n15202));
    defparam n15199_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15967_bdd_4_lut (.I0(n15967), .I1(\REG.mem_21_25 ), .I2(\REG.mem_20_25 ), 
            .I3(rd_addr_r[1]), .O(n13662));
    defparam n15967_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i572_573 (.Q(\REG.mem_5_18 ), .C(FIFO_CLK_c), .D(n5776));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5026_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_28_6 ), .O(n6500));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5026_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i569_570 (.Q(\REG.mem_5_17 ), .C(FIFO_CLK_c), .D(n5775));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5025_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_28_5 ), .O(n6499));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5025_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i566_567 (.Q(\REG.mem_5_16 ), .C(FIFO_CLK_c), .D(n5774));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5024_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_28_4 ), .O(n6498));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5024_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i563_564 (.Q(\REG.mem_5_15 ), .C(FIFO_CLK_c), .D(n5773));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13606 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_25 ), 
            .I2(\REG.mem_15_25 ), .I3(rd_addr_r[1]), .O(n15961));
    defparam rd_addr_r_0__bdd_4_lut_13606.LUT_INIT = 16'he4aa;
    SB_LUT4 i5023_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_28_3 ), .O(n6497));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5023_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5129_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_31_13 ), .O(n6603));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5129_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5128_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_31_12 ), .O(n6602));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5128_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5127_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_31_11 ), .O(n6601));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5127_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5126_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_31_10 ), .O(n6600));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5126_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i560_561 (.Q(\REG.mem_5_14 ), .C(FIFO_CLK_c), .D(n5772));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5125_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_31_9 ), .O(n6599));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5125_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5124_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_31_8 ), .O(n6598));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5124_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15961_bdd_4_lut (.I0(n15961), .I1(\REG.mem_13_25 ), .I2(\REG.mem_12_25 ), 
            .I3(rd_addr_r[1]), .O(n13668));
    defparam n15961_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5022_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_28_2 ), .O(n6496));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5022_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5123_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_31_7 ), .O(n6597));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5123_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5122_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_31_6 ), .O(n6596));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5122_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4156_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_0_18 ), .O(n5630));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4156_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13601 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_20 ), 
            .I2(\REG.mem_31_20 ), .I3(rd_addr_r[1]), .O(n15955));
    defparam rd_addr_r_0__bdd_4_lut_13601.LUT_INIT = 16'he4aa;
    SB_LUT4 n15955_bdd_4_lut (.I0(n15955), .I1(\REG.mem_29_20 ), .I2(\REG.mem_28_20 ), 
            .I3(rd_addr_r[1]), .O(n14235));
    defparam n15955_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12966 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_24 ), 
            .I2(\REG.mem_23_24 ), .I3(rd_addr_r[1]), .O(n15187));
    defparam rd_addr_r_0__bdd_4_lut_12966.LUT_INIT = 16'he4aa;
    SB_LUT4 n15187_bdd_4_lut (.I0(n15187), .I1(\REG.mem_21_24 ), .I2(\REG.mem_20_24 ), 
            .I3(rd_addr_r[1]), .O(n13983));
    defparam n15187_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i557_558 (.Q(\REG.mem_5_13 ), .C(FIFO_CLK_c), .D(n5771));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5021_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_28_1 ), .O(n6495));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5021_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5121_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_31_5 ), .O(n6595));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5121_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5120_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_31_4 ), .O(n6594));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5120_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5119_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_31_3 ), .O(n6593));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5119_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i554_555 (.Q(\REG.mem_5_12 ), .C(FIFO_CLK_c), .D(n5770));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13651 (.I0(rd_addr_r[1]), .I1(n13234), 
            .I2(n13235), .I3(rd_addr_r[2]), .O(n15949));
    defparam rd_addr_r_1__bdd_4_lut_13651.LUT_INIT = 16'he4aa;
    SB_LUT4 n15949_bdd_4_lut (.I0(n15949), .I1(n13232), .I2(n13231), .I3(rd_addr_r[2]), 
            .O(n13268));
    defparam n15949_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12956 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_12 ), 
            .I2(\REG.mem_15_12 ), .I3(rd_addr_r[1]), .O(n15181));
    defparam rd_addr_r_0__bdd_4_lut_12956.LUT_INIT = 16'he4aa;
    SB_LUT4 i5118_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_31_2 ), .O(n6592));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5118_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i551_552 (.Q(\REG.mem_5_11 ), .C(FIFO_CLK_c), .D(n5769));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5117_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_31_1 ), .O(n6591));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5117_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12077_3_lut (.I0(\REG.mem_24_3 ), .I1(\REG.mem_25_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14188));
    defparam i12077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n15181_bdd_4_lut (.I0(n15181), .I1(\REG.mem_13_12 ), .I2(\REG.mem_12_12 ), 
            .I3(rd_addr_r[1]), .O(n15184));
    defparam n15181_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13596 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_25 ), 
            .I2(\REG.mem_3_25 ), .I3(rd_addr_r[1]), .O(n15943));
    defparam rd_addr_r_0__bdd_4_lut_13596.LUT_INIT = 16'he4aa;
    SB_LUT4 n15943_bdd_4_lut (.I0(n15943), .I1(\REG.mem_1_25 ), .I2(\REG.mem_0_25 ), 
            .I3(rd_addr_r[1]), .O(n13683));
    defparam n15943_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i548_549 (.Q(\REG.mem_5_10 ), .C(FIFO_CLK_c), .D(n5768));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5116_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_31_0 ), .O(n6590));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5116_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12078_3_lut (.I0(\REG.mem_26_3 ), .I1(\REG.mem_27_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14189));
    defparam i12078_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i545_546 (.Q(\REG.mem_5_9 ), .C(FIFO_CLK_c), .D(n5767));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i12084_3_lut (.I0(\REG.mem_30_3 ), .I1(\REG.mem_31_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14195));
    defparam i12084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i34_2_lut_3_lut (.I0(n10_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n34));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i34_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i542_543 (.Q(\REG.mem_5_8 ), .C(FIFO_CLK_c), .D(n5766));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i12083_3_lut (.I0(\REG.mem_28_3 ), .I1(\REG.mem_29_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14194));
    defparam i12083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5020_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_28_0 ), .O(n6494));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5020_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13591 (.I0(rd_addr_r[1]), .I1(n13594), 
            .I2(n13595), .I3(rd_addr_r[2]), .O(n15937));
    defparam rd_addr_r_1__bdd_4_lut_13591.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12951 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_6 ), 
            .I2(\REG.mem_27_6 ), .I3(rd_addr_r[1]), .O(n15175));
    defparam rd_addr_r_0__bdd_4_lut_12951.LUT_INIT = 16'he4aa;
    SB_LUT4 n15937_bdd_4_lut (.I0(n15937), .I1(n13562), .I2(n13561), .I3(rd_addr_r[2]), 
            .O(n13691));
    defparam n15937_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i539_540 (.Q(\REG.mem_5_7 ), .C(FIFO_CLK_c), .D(n5765));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4157_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_0_7 ), .O(n5631));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4157_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15175_bdd_4_lut (.I0(n15175), .I1(\REG.mem_25_6 ), .I2(\REG.mem_24_6 ), 
            .I3(rd_addr_r[1]), .O(n13986));
    defparam n15175_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i50_2_lut_3_lut_4_lut (.I0(n10_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n10));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i50_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13581 (.I0(rd_addr_r[1]), .I1(n13255), 
            .I2(n13256), .I3(rd_addr_r[2]), .O(n15931));
    defparam rd_addr_r_1__bdd_4_lut_13581.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12946 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_24 ), 
            .I2(\REG.mem_27_24 ), .I3(rd_addr_r[1]), .O(n15169));
    defparam rd_addr_r_0__bdd_4_lut_12946.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i51_2_lut_3_lut_4_lut (.I0(n10_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n26));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i51_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_DFF i146_147 (.Q(\REG.mem_1_4 ), .C(FIFO_CLK_c), .D(n5596));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4159_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_0_16 ), .O(n5633));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4159_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i536_537 (.Q(\REG.mem_5_6 ), .C(FIFO_CLK_c), .D(n5764));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n15169_bdd_4_lut (.I0(n15169), .I1(\REG.mem_25_24 ), .I2(\REG.mem_24_24 ), 
            .I3(rd_addr_r[1]), .O(n13989));
    defparam n15169_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15931_bdd_4_lut (.I0(n15931), .I1(n13250), .I2(n13249), .I3(rd_addr_r[2]), 
            .O(n13280));
    defparam n15931_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i149_150 (.Q(\REG.mem_1_5 ), .C(FIFO_CLK_c), .D(n5595));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13021 (.I0(rd_addr_r[1]), .I1(n14215), 
            .I2(n14216), .I3(rd_addr_r[2]), .O(n15163));
    defparam rd_addr_r_1__bdd_4_lut_13021.LUT_INIT = 16'he4aa;
    SB_LUT4 n15163_bdd_4_lut (.I0(n15163), .I1(n14213), .I2(n14212), .I3(rd_addr_r[2]), 
            .O(n15166));
    defparam n15163_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i152_153 (.Q(\REG.mem_1_6 ), .C(FIFO_CLK_c), .D(n5594));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4155_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_0_19 ), .O(n5629));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4155_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i155_156 (.Q(\REG.mem_1_7 ), .C(FIFO_CLK_c), .D(n5593));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12941 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_6 ), 
            .I2(\REG.mem_31_6 ), .I3(rd_addr_r[1]), .O(n15151));
    defparam rd_addr_r_0__bdd_4_lut_12941.LUT_INIT = 16'he4aa;
    SB_LUT4 i4635_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_15_31 ), .O(n6109));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4635_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut (.I0(rd_addr_r[3]), .I1(n14158), .I2(n14159), 
            .I3(rd_addr_r[4]), .O(n15913));
    defparam rd_addr_r_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n15913_bdd_4_lut (.I0(n15913), .I1(n14141), .I2(n14140), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[23]));
    defparam n15913_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4634_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_15_30 ), .O(n6108));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4634_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4539_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_12_31 ), .O(n6013));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4539_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4633_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_15_29 ), .O(n6107));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4633_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13576 (.I0(rd_addr_r[1]), .I1(n13696), 
            .I2(n13697), .I3(rd_addr_r[2]), .O(n15907));
    defparam rd_addr_r_1__bdd_4_lut_13576.LUT_INIT = 16'he4aa;
    SB_LUT4 n15907_bdd_4_lut (.I0(n15907), .I1(n13643), .I2(n13642), .I3(rd_addr_r[2]), 
            .O(n13706));
    defparam n15907_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4538_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_12_30 ), .O(n6012));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4538_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4632_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_15_28 ), .O(n6106));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4632_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4537_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_12_29 ), .O(n6011));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4537_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i224_225 (.Q(\REG.mem_1_30 ), .C(FIFO_CLK_c), .D(n5590));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4631_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_15_27 ), .O(n6105));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4631_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4630_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_15_26 ), .O(n6104));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4630_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4629_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_15_25 ), .O(n6103));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4629_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_13561 (.I0(rd_addr_r[3]), .I1(n13567), 
            .I2(n13568), .I3(rd_addr_r[4]), .O(n15901));
    defparam rd_addr_r_3__bdd_4_lut_13561.LUT_INIT = 16'he4aa;
    SB_LUT4 n14491_bdd_4_lut (.I0(n14491), .I1(\REG.mem_21_12 ), .I2(\REG.mem_20_12 ), 
            .I3(rd_addr_r[1]), .O(n14494));
    defparam n14491_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15901_bdd_4_lut (.I0(n15901), .I1(n14129), .I2(n14128), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[4]));
    defparam n15901_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15151_bdd_4_lut (.I0(n15151), .I1(\REG.mem_29_6 ), .I2(\REG.mem_28_6 ), 
            .I3(rd_addr_r[1]), .O(n13995));
    defparam n15151_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4628_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_15_24 ), .O(n6102));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4628_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4627_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_15_23 ), .O(n6101));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4627_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12926 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_8 ), 
            .I2(\REG.mem_31_8 ), .I3(rd_addr_r[1]), .O(n15145));
    defparam rd_addr_r_0__bdd_4_lut_12926.LUT_INIT = 16'he4aa;
    SB_LUT4 i4536_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_12_28 ), .O(n6010));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4536_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4626_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_15_22 ), .O(n6100));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4626_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15145_bdd_4_lut (.I0(n15145), .I1(\REG.mem_29_8 ), .I2(\REG.mem_28_8 ), 
            .I3(rd_addr_r[1]), .O(n13998));
    defparam n15145_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4625_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_15_21 ), .O(n6099));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4625_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13556 (.I0(rd_addr_r[1]), .I1(n13261), 
            .I2(n13262), .I3(rd_addr_r[2]), .O(n15895));
    defparam rd_addr_r_1__bdd_4_lut_13556.LUT_INIT = 16'he4aa;
    SB_LUT4 i4624_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_15_20 ), .O(n6098));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4624_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4623_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_15_19 ), .O(n6097));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4623_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15895_bdd_4_lut (.I0(n15895), .I1(n13253), .I2(n13252), .I3(rd_addr_r[2]), 
            .O(n13304));
    defparam n15895_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY wp_sync2_r_5__I_0_135_add_2_2 (.CI(VCC_net), .I0(wp_sync_w[0]), 
            .I1(n1[0]), .CO(n12066));
    SB_LUT4 i4535_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_12_27 ), .O(n6009));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4535_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4622_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_15_18 ), .O(n6096));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4622_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_13031 (.I0(rd_addr_r[3]), .I1(n15022), 
            .I2(n13454), .I3(rd_addr_r[4]), .O(n15139));
    defparam rd_addr_r_3__bdd_4_lut_13031.LUT_INIT = 16'he4aa;
    SB_DFF i218_219 (.Q(\REG.mem_1_28 ), .C(FIFO_CLK_c), .D(n5589));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4621_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_15_17 ), .O(n6095));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4621_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4534_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_12_26 ), .O(n6008));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4534_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4620_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_15_16 ), .O(n6094));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4620_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF wp_sync2_r__i0 (.Q(wp_sync2_r[0]), .C(SLM_CLK_c), .D(n5588));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_LUT4 i4619_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_15_15 ), .O(n6093));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4619_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i191_192 (.Q(\REG.mem_1_19 ), .C(FIFO_CLK_c), .D(n5587));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i533_534 (.Q(\REG.mem_5_5 ), .C(FIFO_CLK_c), .D(n5763));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4533_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_12_25 ), .O(n6007));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4533_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15139_bdd_4_lut (.I0(n15139), .I1(n13838), .I2(n13837), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[17]));
    defparam n15139_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12448 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_26 ), 
            .I2(\REG.mem_7_26 ), .I3(rd_addr_r[1]), .O(n14563));
    defparam rd_addr_r_0__bdd_4_lut_12448.LUT_INIT = 16'he4aa;
    SB_LUT4 i4532_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_12_24 ), .O(n6006));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4532_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14563_bdd_4_lut (.I0(n14563), .I1(\REG.mem_5_26 ), .I2(\REG.mem_4_26 ), 
            .I3(rd_addr_r[1]), .O(n14566));
    defparam n14563_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4531_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_12_23 ), .O(n6005));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4531_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i530_531 (.Q(\REG.mem_5_4 ), .C(FIFO_CLK_c), .D(n5762));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4160_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_0_15 ), .O(n5634));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4160_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13546 (.I0(rd_addr_r[1]), .I1(n13201), 
            .I2(n13202), .I3(rd_addr_r[2]), .O(n15889));
    defparam rd_addr_r_1__bdd_4_lut_13546.LUT_INIT = 16'he4aa;
    SB_DFF i527_528 (.Q(\REG.mem_5_3 ), .C(FIFO_CLK_c), .D(n5761));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4163_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_0_14 ), .O(n5637));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4163_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15889_bdd_4_lut (.I0(n15889), .I1(n13199), .I2(n13198), .I3(rd_addr_r[2]), 
            .O(n13963));
    defparam n15889_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4618_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_15_14 ), .O(n6092));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4618_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4617_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_15_13 ), .O(n6091));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4617_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i524_525 (.Q(\REG.mem_5_2 ), .C(FIFO_CLK_c), .D(n5760));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i521_522 (.Q(\REG.mem_5_1 ), .C(FIFO_CLK_c), .D(n5759));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13541 (.I0(rd_addr_r[1]), .I1(n13111), 
            .I2(n13112), .I3(rd_addr_r[2]), .O(n15883));
    defparam rd_addr_r_1__bdd_4_lut_13541.LUT_INIT = 16'he4aa;
    SB_LUT4 i4616_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_15_12 ), .O(n6090));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4616_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4615_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_15_11 ), .O(n6089));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4615_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12513 (.I0(rd_addr_r[2]), .I1(n14232), 
            .I2(n14235), .I3(rd_addr_r[3]), .O(n14557));
    defparam rd_addr_r_2__bdd_4_lut_12513.LUT_INIT = 16'he4aa;
    SB_LUT4 i4614_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_15_10 ), .O(n6088));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4614_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4613_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_15_9 ), .O(n6087));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4613_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4612_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_15_8 ), .O(n6086));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4612_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4530_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_12_22 ), .O(n6004));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4530_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4611_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_15_7 ), .O(n6085));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4611_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4610_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_15_6 ), .O(n6084));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4610_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15883_bdd_4_lut (.I0(n15883), .I1(n13106), .I2(n13105), .I3(rd_addr_r[2]), 
            .O(n13124));
    defparam n15883_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4609_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_15_5 ), .O(n6083));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4609_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF wp_sync1_r__i0 (.Q(wp_sync1_r[0]), .C(SLM_CLK_c), .D(n5586));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF i518_519 (.Q(\REG.mem_5_0 ), .C(FIFO_CLK_c), .D(n5758));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4608_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_15_4 ), .O(n6082));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4608_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i515_516 (.Q(\REG.mem_4_31 ), .C(FIFO_CLK_c), .D(n5757));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4607_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_15_3 ), .O(n6081));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4607_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i512_513 (.Q(\REG.mem_4_30 ), .C(FIFO_CLK_c), .D(n5756));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4529_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_12_21 ), .O(n6003));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4529_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4606_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_15_2 ), .O(n6080));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4606_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4528_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_12_20 ), .O(n6002));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4528_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4605_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_15_1 ), .O(n6079));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4605_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4527_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_12_19 ), .O(n6001));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4527_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13536 (.I0(rd_addr_r[1]), .I1(n13624), 
            .I2(n13625), .I3(rd_addr_r[2]), .O(n15877));
    defparam rd_addr_r_1__bdd_4_lut_13536.LUT_INIT = 16'he4aa;
    SB_LUT4 i4604_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_15_0 ), .O(n6078));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4604_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5115_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_30_31 ), .O(n6589));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5115_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15877_bdd_4_lut (.I0(n15877), .I1(n13592), .I2(n13591), .I3(rd_addr_r[2]), 
            .O(n13730));
    defparam n15877_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4164_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_0_13 ), .O(n5638));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4164_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13531 (.I0(rd_addr_r[1]), .I1(n13285), 
            .I2(n13286), .I3(rd_addr_r[2]), .O(n15871));
    defparam rd_addr_r_1__bdd_4_lut_13531.LUT_INIT = 16'he4aa;
    SB_LUT4 i5114_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_30_30 ), .O(n6588));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5114_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i509_510 (.Q(\REG.mem_4_29 ), .C(FIFO_CLK_c), .D(n5755));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n15871_bdd_4_lut (.I0(n15871), .I1(n13283), .I2(n13282), .I3(rd_addr_r[2]), 
            .O(n13316));
    defparam n15871_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12921 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_0 ), 
            .I2(\REG.mem_15_0 ), .I3(rd_addr_r[1]), .O(n15127));
    defparam rd_addr_r_0__bdd_4_lut_12921.LUT_INIT = 16'he4aa;
    SB_LUT4 n15127_bdd_4_lut (.I0(n15127), .I1(\REG.mem_13_0 ), .I2(\REG.mem_12_0 ), 
            .I3(rd_addr_r[1]), .O(n13479));
    defparam n15127_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5113_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_30_29 ), .O(n6587));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5113_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13526 (.I0(rd_addr_r[1]), .I1(n13657), 
            .I2(n13658), .I3(rd_addr_r[2]), .O(n15865));
    defparam rd_addr_r_1__bdd_4_lut_13526.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_r_5__I_0_123_i5_3_lut (.I0(wr_addr_r[4]), .I1(wr_addr_p1_w[4]), 
            .I2(wr_fifo_en_w), .I3(GND_net), .O(\wr_addr_nxt_c[4] ));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_5__I_0_123_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i506_507 (.Q(\REG.mem_4_28 ), .C(FIFO_CLK_c), .D(n5754));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i503_504 (.Q(\REG.mem_4_27 ), .C(FIFO_CLK_c), .D(n5753));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i500_501 (.Q(\REG.mem_4_26 ), .C(FIFO_CLK_c), .D(n5752));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i497_498 (.Q(\REG.mem_4_25 ), .C(FIFO_CLK_c), .D(n5751));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i494_495 (.Q(\REG.mem_4_24 ), .C(FIFO_CLK_c), .D(n5750));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i491_492 (.Q(\REG.mem_4_23 ), .C(FIFO_CLK_c), .D(n5749));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i488_489 (.Q(\REG.mem_4_22 ), .C(FIFO_CLK_c), .D(n5748));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i485_486 (.Q(\REG.mem_4_21 ), .C(FIFO_CLK_c), .D(n5747));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i221_222 (.Q(\REG.mem_1_29 ), .C(FIFO_CLK_c), .D(n5585));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rd_addr_r__i0 (.Q(rd_addr_r[0]), .C(SLM_CLK_c), .D(n5584));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF i206_207 (.Q(\REG.mem_1_24 ), .C(FIFO_CLK_c), .D(n5583));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync2_r__i0 (.Q(rp_sync2_r[0]), .C(FIFO_CLK_c), .D(n5582));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF i158_159 (.Q(\REG.mem_1_8 ), .C(FIFO_CLK_c), .D(n5581));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync1_r__i0 (.Q(rp_sync1_r[0]), .C(FIFO_CLK_c), .D(n5580));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF i62_63 (.Q(\REG.mem_0_8 ), .C(FIFO_CLK_c), .D(n5579));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i161_162 (.Q(\REG.mem_1_9 ), .C(FIFO_CLK_c), .D(n5577));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i482_483 (.Q(\REG.mem_4_20 ), .C(FIFO_CLK_c), .D(n5746));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14557_bdd_4_lut (.I0(n14557), .I1(n14229), .I2(n14226), .I3(rd_addr_r[3]), 
            .O(n14560));
    defparam n14557_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4165_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_0_12 ), .O(n5639));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4165_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4526_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_12_18 ), .O(n6000));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4526_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5112_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_30_28 ), .O(n6586));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5112_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5111_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_30_27 ), .O(n6585));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5111_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i479_480 (.Q(\REG.mem_4_19 ), .C(FIFO_CLK_c), .D(n5745));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i476_477 (.Q(\REG.mem_4_18 ), .C(FIFO_CLK_c), .D(n5744));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i473_474 (.Q(\REG.mem_4_17 ), .C(FIFO_CLK_c), .D(n5743));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i470_471 (.Q(\REG.mem_4_16 ), .C(FIFO_CLK_c), .D(n5742));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i467_468 (.Q(\REG.mem_4_15 ), .C(FIFO_CLK_c), .D(n5741));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i464_465 (.Q(\REG.mem_4_14 ), .C(FIFO_CLK_c), .D(n5740));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i461_462 (.Q(\REG.mem_4_13 ), .C(FIFO_CLK_c), .D(n5739));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i458_459 (.Q(\REG.mem_4_12 ), .C(FIFO_CLK_c), .D(n5738));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i164_165 (.Q(\REG.mem_1_10 ), .C(FIFO_CLK_c), .D(n5574));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i227_228 (.Q(\REG.mem_1_31 ), .C(FIFO_CLK_c), .D(n5572));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i167_168 (.Q(\REG.mem_1_11 ), .C(FIFO_CLK_c), .D(n5571));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i41_42 (.Q(\REG.mem_0_1 ), .C(FIFO_CLK_c), .D(n5570));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i44_45 (.Q(\REG.mem_0_2 ), .C(FIFO_CLK_c), .D(n5569));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i53_54 (.Q(\REG.mem_0_5 ), .C(FIFO_CLK_c), .D(n5568));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i455_456 (.Q(\REG.mem_4_11 ), .C(FIFO_CLK_c), .D(n5737));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n15865_bdd_4_lut (.I0(n15865), .I1(n13616), .I2(n13615), .I3(rd_addr_r[2]), 
            .O(n13742));
    defparam n15865_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5110_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_30_26 ), .O(n6584));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5110_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i452_453 (.Q(\REG.mem_4_10 ), .C(FIFO_CLK_c), .D(n5736));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i449_450 (.Q(\REG.mem_4_9 ), .C(FIFO_CLK_c), .D(n5735));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i446_447 (.Q(\REG.mem_4_8 ), .C(FIFO_CLK_c), .D(n5734));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i443_444 (.Q(\REG.mem_4_7 ), .C(FIFO_CLK_c), .D(n5733));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i440_441 (.Q(\REG.mem_4_6 ), .C(FIFO_CLK_c), .D(n5732));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i437_438 (.Q(\REG.mem_4_5 ), .C(FIFO_CLK_c), .D(n5731));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i434_435 (.Q(\REG.mem_4_4 ), .C(FIFO_CLK_c), .D(n5730));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i431_432 (.Q(\REG.mem_4_3 ), .C(FIFO_CLK_c), .D(n5729));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i185_186 (.Q(\REG.mem_1_17 ), .C(FIFO_CLK_c), .D(n5567));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i194_195 (.Q(\REG.mem_1_20 ), .C(FIFO_CLK_c), .D(n5565));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i170_171 (.Q(\REG.mem_1_12 ), .C(FIFO_CLK_c), .D(n5564));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i47_48 (.Q(\REG.mem_0_3 ), .C(FIFO_CLK_c), .D(n5563));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i50_51 (.Q(\REG.mem_0_4 ), .C(FIFO_CLK_c), .D(n5562));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i56_57 (.Q(\REG.mem_0_6 ), .C(FIFO_CLK_c), .D(n5561));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i173_174 (.Q(\REG.mem_1_13 ), .C(FIFO_CLK_c), .D(n5560));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i176_177 (.Q(\REG.mem_1_14 ), .C(FIFO_CLK_c), .D(n5559));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i179_180 (.Q(\REG.mem_1_15 ), .C(FIFO_CLK_c), .D(n5558));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5109_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_30_25 ), .O(n6583));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5109_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5108_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_30_24 ), .O(n6582));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5108_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4525_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_12_17 ), .O(n5999));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4525_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i182_183 (.Q(\REG.mem_1_16 ), .C(FIFO_CLK_c), .D(n5557));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5107_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_30_23 ), .O(n6581));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5107_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4524_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_12_16 ), .O(n5998));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4524_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i209_210 (.Q(\REG.mem_1_25 ), .C(FIFO_CLK_c), .D(n5556));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5106_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_30_22 ), .O(n6580));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5106_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13586 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_10 ), 
            .I2(\REG.mem_27_10 ), .I3(rd_addr_r[1]), .O(n15859));
    defparam rd_addr_r_0__bdd_4_lut_13586.LUT_INIT = 16'he4aa;
    SB_LUT4 i4523_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_12_15 ), .O(n5997));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4523_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15859_bdd_4_lut (.I0(n15859), .I1(\REG.mem_25_10 ), .I2(\REG.mem_24_10 ), 
            .I3(rd_addr_r[1]), .O(n15862));
    defparam n15859_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4522_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_12_14 ), .O(n5996));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4522_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i197_198 (.Q(\REG.mem_1_21 ), .C(FIFO_CLK_c), .D(n5555));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4763_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_19_31 ), .O(n6237));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4763_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_r_5__I_0_123_i3_3_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_w[2]), 
            .I2(wr_fifo_en_w), .I3(GND_net), .O(\wr_addr_nxt_c[2] ));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_5__I_0_123_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4762_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_19_30 ), .O(n6236));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4762_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF wr_addr_r__i0 (.Q(\wr_addr_r[0] ), .C(FIFO_CLK_c), .D(n5554));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 i4761_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_19_29 ), .O(n6235));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4761_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5105_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_30_21 ), .O(n6579));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5105_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4760_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_19_28 ), .O(n6234));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4760_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4759_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_19_27 ), .O(n6233));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4759_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5104_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_30_20 ), .O(n6578));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5104_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5103_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_30_19 ), .O(n6577));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5103_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i212_213 (.Q(\REG.mem_1_26 ), .C(FIFO_CLK_c), .D(n5551));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5102_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_30_18 ), .O(n6576));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5102_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i200_201 (.Q(\REG.mem_1_22 ), .C(FIFO_CLK_c), .D(n5550));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5101_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_30_17 ), .O(n6575));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5101_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i428_429 (.Q(\REG.mem_4_2 ), .C(FIFO_CLK_c), .D(n5728));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i425_426 (.Q(\REG.mem_4_1 ), .C(FIFO_CLK_c), .D(n5727));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i422_423 (.Q(\REG.mem_4_0 ), .C(FIFO_CLK_c), .D(n5726));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4758_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_19_26 ), .O(n6232));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4758_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i419_420 (.Q(\REG.mem_3_31 ), .C(FIFO_CLK_c), .D(n5725));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i416_417 (.Q(\REG.mem_3_30 ), .C(FIFO_CLK_c), .D(n5724));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i413_414 (.Q(\REG.mem_3_29 ), .C(FIFO_CLK_c), .D(n5723));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12907 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_28 ), 
            .I2(\REG.mem_31_28 ), .I3(rd_addr_r[1]), .O(n15115));
    defparam rd_addr_r_0__bdd_4_lut_12907.LUT_INIT = 16'he4aa;
    SB_DFF i410_411 (.Q(\REG.mem_3_28 ), .C(FIFO_CLK_c), .D(n5722));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4757_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_19_25 ), .O(n6231));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4757_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i407_408 (.Q(\REG.mem_3_27 ), .C(FIFO_CLK_c), .D(n5721));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i404_405 (.Q(\REG.mem_3_26 ), .C(FIFO_CLK_c), .D(n5720));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i401_402 (.Q(\REG.mem_3_25 ), .C(FIFO_CLK_c), .D(n5719));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i398_399 (.Q(\REG.mem_3_24 ), .C(FIFO_CLK_c), .D(n5718));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4756_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_19_24 ), .O(n6230));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4756_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i395_396 (.Q(\REG.mem_3_23 ), .C(FIFO_CLK_c), .D(n5717));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i392_393 (.Q(\REG.mem_3_22 ), .C(FIFO_CLK_c), .D(n5716));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i389_390 (.Q(\REG.mem_3_21 ), .C(FIFO_CLK_c), .D(n5715));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i386_387 (.Q(\REG.mem_3_20 ), .C(FIFO_CLK_c), .D(n5714));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4521_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_12_13 ), .O(n5995));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4521_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4755_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_19_23 ), .O(n6229));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4755_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4520_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_12_12 ), .O(n5994));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4520_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4754_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_19_22 ), .O(n6228));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4754_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4753_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_19_21 ), .O(n6227));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4753_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i383_384 (.Q(\REG.mem_3_19 ), .C(FIFO_CLK_c), .D(n5713));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i380_381 (.Q(\REG.mem_3_18 ), .C(FIFO_CLK_c), .D(n5712));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5100_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_30_16 ), .O(n6574));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5100_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4752_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_19_20 ), .O(n6226));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4752_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4751_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_19_19 ), .O(n6225));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4751_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15115_bdd_4_lut (.I0(n15115), .I1(\REG.mem_29_28 ), .I2(\REG.mem_28_28 ), 
            .I3(rd_addr_r[1]), .O(n14004));
    defparam n15115_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5099_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_30_15 ), .O(n6573));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5099_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4750_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_19_18 ), .O(n6224));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4750_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i377_378 (.Q(\REG.mem_3_17 ), .C(FIFO_CLK_c), .D(n5711));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13521 (.I0(rd_addr_r[1]), .I1(n13300), 
            .I2(n13301), .I3(rd_addr_r[2]), .O(n15847));
    defparam rd_addr_r_1__bdd_4_lut_13521.LUT_INIT = 16'he4aa;
    SB_LUT4 i4749_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_19_17 ), .O(n6223));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4749_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12897 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_5 ), 
            .I2(\REG.mem_3_5 ), .I3(rd_addr_r[1]), .O(n15109));
    defparam rd_addr_r_0__bdd_4_lut_12897.LUT_INIT = 16'he4aa;
    SB_DFF i374_375 (.Q(\REG.mem_3_16 ), .C(FIFO_CLK_c), .D(n5710));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4748_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_19_16 ), .O(n6222));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4748_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i371_372 (.Q(\REG.mem_3_15 ), .C(FIFO_CLK_c), .D(n5709));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4127_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_0_0 ), .O(n5601));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4127_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5098_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_30_14 ), .O(n6572));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5098_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5097_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_30_13 ), .O(n6571));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5097_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4167_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_0_11 ), .O(n5641));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4167_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4747_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_19_15 ), .O(n6221));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4747_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i368_369 (.Q(\REG.mem_3_14 ), .C(FIFO_CLK_c), .D(n5708));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4168_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_0_10 ), .O(n5642));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4168_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4105_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_0_8 ), .O(n5579));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4105_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4158_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_0_17 ), .O(n5632));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4158_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i365_366 (.Q(\REG.mem_3_13 ), .C(FIFO_CLK_c), .D(n5707));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5096_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_30_12 ), .O(n6570));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5096_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4089_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_0_3 ), .O(n5563));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4089_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4746_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_19_14 ), .O(n6220));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4746_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i362_363 (.Q(\REG.mem_3_12 ), .C(FIFO_CLK_c), .D(n5706));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5095_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_30_11 ), .O(n6569));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5095_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15847_bdd_4_lut (.I0(n15847), .I1(n13298), .I2(n13297), .I3(rd_addr_r[2]), 
            .O(n13325));
    defparam n15847_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i359_360 (.Q(\REG.mem_3_11 ), .C(FIFO_CLK_c), .D(n5705));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5094_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_30_10 ), .O(n6568));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5094_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13506 (.I0(rd_addr_r[1]), .I1(n13264), 
            .I2(n13265), .I3(rd_addr_r[2]), .O(n15841));
    defparam rd_addr_r_1__bdd_4_lut_13506.LUT_INIT = 16'he4aa;
    SB_LUT4 i4745_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_19_13 ), .O(n6219));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4745_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15109_bdd_4_lut (.I0(n15109), .I1(\REG.mem_1_5 ), .I2(\REG.mem_0_5 ), 
            .I3(rd_addr_r[1]), .O(n14007));
    defparam n15109_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4744_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_19_12 ), .O(n6218));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4744_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5093_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_30_9 ), .O(n6567));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5093_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4743_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_19_11 ), .O(n6217));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4743_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5092_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_30_8 ), .O(n6566));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5092_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12438 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_4 ), 
            .I2(\REG.mem_15_4 ), .I3(rd_addr_r[1]), .O(n14551));
    defparam rd_addr_r_0__bdd_4_lut_12438.LUT_INIT = 16'he4aa;
    SB_LUT4 i5091_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_30_7 ), .O(n6565));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5091_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4742_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_19_10 ), .O(n6216));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4742_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15841_bdd_4_lut (.I0(n15841), .I1(n13259), .I2(n13258), .I3(rd_addr_r[2]), 
            .O(n13891));
    defparam n15841_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4741_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_19_9 ), .O(n6215));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4741_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4519_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_12_11 ), .O(n5993));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4519_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5090_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_30_6 ), .O(n6564));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5090_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5089_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_30_5 ), .O(n6563));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5089_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5088_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_30_4 ), .O(n6562));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5088_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4518_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_12_10 ), .O(n5992));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4518_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5087_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_30_3 ), .O(n6561));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5087_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4740_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_19_8 ), .O(n6214));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4740_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12936 (.I0(rd_addr_r[1]), .I1(n13375), 
            .I2(n13376), .I3(rd_addr_r[2]), .O(n15103));
    defparam rd_addr_r_1__bdd_4_lut_12936.LUT_INIT = 16'he4aa;
    SB_LUT4 i5086_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_30_2 ), .O(n6560));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5086_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4739_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_19_7 ), .O(n6213));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4739_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14551_bdd_4_lut (.I0(n14551), .I1(\REG.mem_13_4 ), .I2(\REG.mem_12_4 ), 
            .I3(rd_addr_r[1]), .O(n14554));
    defparam n14551_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4738_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_19_6 ), .O(n6212));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4738_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15103_bdd_4_lut (.I0(n15103), .I1(n13370), .I2(n13369), .I3(rd_addr_r[2]), 
            .O(n13484));
    defparam n15103_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4737_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_19_5 ), .O(n6211));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4737_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5085_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_30_1 ), .O(n6559));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5085_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5084_3_lut_4_lut (.I0(n32_adj_1376), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_30_0 ), .O(n6558));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5084_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4517_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_12_9 ), .O(n5991));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4517_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13516 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_25 ), 
            .I2(\REG.mem_7_25 ), .I3(rd_addr_r[1]), .O(n15829));
    defparam rd_addr_r_0__bdd_4_lut_13516.LUT_INIT = 16'he4aa;
    SB_LUT4 i4736_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_19_4 ), .O(n6210));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4736_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15829_bdd_4_lut (.I0(n15829), .I1(\REG.mem_5_25 ), .I2(\REG.mem_4_25 ), 
            .I3(rd_addr_r[1]), .O(n13761));
    defparam n15829_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4735_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_19_3 ), .O(n6209));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4735_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i32_2_lut_3_lut (.I0(n8_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n32_adj_1376));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i32_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12887 (.I0(rd_addr_r[1]), .I1(n13861), 
            .I2(n13862), .I3(rd_addr_r[2]), .O(n15097));
    defparam rd_addr_r_1__bdd_4_lut_12887.LUT_INIT = 16'he4aa;
    SB_LUT4 i4516_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_12_8 ), .O(n5990));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4516_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13491 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_25 ), 
            .I2(\REG.mem_11_25 ), .I3(rd_addr_r[1]), .O(n15823));
    defparam rd_addr_r_0__bdd_4_lut_13491.LUT_INIT = 16'he4aa;
    SB_LUT4 i4734_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_19_2 ), .O(n6208));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4734_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10952_3_lut (.I0(\REG.mem_0_11 ), .I1(\REG.mem_1_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13063));
    defparam i10952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n15823_bdd_4_lut (.I0(n15823), .I1(\REG.mem_9_25 ), .I2(\REG.mem_8_25 ), 
            .I3(rd_addr_r[1]), .O(n13764));
    defparam n15823_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10953_3_lut (.I0(\REG.mem_2_11 ), .I1(\REG.mem_3_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13064));
    defparam i10953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4733_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_19_1 ), .O(n6207));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4733_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4732_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_19_0 ), .O(n6206));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4732_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4515_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_12_7 ), .O(n5989));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4515_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_addr_nxt_c_5__I_0_136_i4_2_lut_4_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_w[3]), 
            .I2(wr_fifo_en_w), .I3(\wr_addr_nxt_c[4] ), .O(wr_grey_w[3]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_5__I_0_136_i4_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 n15097_bdd_4_lut (.I0(n15097), .I1(n13118), .I2(n13117), .I3(rd_addr_r[2]), 
            .O(n13154));
    defparam n15097_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13486 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_16 ), 
            .I2(\REG.mem_11_16 ), .I3(rd_addr_r[1]), .O(n15817));
    defparam rd_addr_r_0__bdd_4_lut_13486.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_nxt_c_5__I_0_136_i3_2_lut_4_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_w[3]), 
            .I2(wr_fifo_en_w), .I3(\wr_addr_nxt_c[2] ), .O(wr_grey_w[2]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_5__I_0_136_i3_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4514_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_12_6 ), .O(n5988));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4514_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5455_2_lut_4_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_w[3]), 
            .I2(wr_fifo_en_w), .I3(reset_per_frame), .O(n6929));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i5455_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 n15817_bdd_4_lut (.I0(n15817), .I1(\REG.mem_9_16 ), .I2(\REG.mem_8_16 ), 
            .I3(rd_addr_r[1]), .O(n13767));
    defparam n15817_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12892 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_16 ), 
            .I2(\REG.mem_27_16 ), .I3(rd_addr_r[1]), .O(n15091));
    defparam rd_addr_r_0__bdd_4_lut_12892.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_nxt_c_5__I_0_136_i5_2_lut_4_lut (.I0(\wr_addr_r[5] ), 
            .I1(wr_addr_p1_w[5]), .I2(wr_fifo_en_w), .I3(\wr_addr_nxt_c[4] ), 
            .O(wr_grey_w[4]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_5__I_0_136_i5_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i5453_2_lut_4_lut (.I0(\wr_addr_r[5] ), .I1(wr_addr_p1_w[5]), 
            .I2(wr_fifo_en_w), .I3(reset_per_frame), .O(n6927));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i5453_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 EnabledDecoder_2_i48_2_lut_3_lut_4_lut (.I0(n8_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n11));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i48_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 n15091_bdd_4_lut (.I0(n15091), .I1(\REG.mem_25_16 ), .I2(\REG.mem_24_16 ), 
            .I3(rd_addr_r[1]), .O(n15094));
    defparam n15091_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4731_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_18_31 ), .O(n6205));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4731_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4730_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_18_30 ), .O(n6204));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4730_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4729_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_18_29 ), .O(n6203));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4729_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i49_2_lut_3_lut_4_lut (.I0(n8_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n27));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i49_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i4513_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_12_5 ), .O(n5987));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4513_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13481 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_22 ), 
            .I2(\REG.mem_15_22 ), .I3(rd_addr_r[1]), .O(n15805));
    defparam rd_addr_r_0__bdd_4_lut_13481.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12877 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_5 ), 
            .I2(\REG.mem_7_5 ), .I3(rd_addr_r[1]), .O(n15085));
    defparam rd_addr_r_0__bdd_4_lut_12877.LUT_INIT = 16'he4aa;
    SB_LUT4 i4728_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_18_28 ), .O(n6202));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4728_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4727_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_18_27 ), .O(n6201));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4727_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15805_bdd_4_lut (.I0(n15805), .I1(\REG.mem_13_22 ), .I2(\REG.mem_12_22 ), 
            .I3(rd_addr_r[1]), .O(n15808));
    defparam n15805_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n15085_bdd_4_lut (.I0(n15085), .I1(\REG.mem_5_5 ), .I2(\REG.mem_4_5 ), 
            .I3(rd_addr_r[1]), .O(n14013));
    defparam n15085_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4512_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_12_4 ), .O(n5986));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4512_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4094_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_0_5 ), .O(n5568));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4094_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4726_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_18_26 ), .O(n6200));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4726_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4725_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_18_25 ), .O(n6199));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4725_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4724_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_18_24 ), .O(n6198));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4724_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4723_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_18_23 ), .O(n6197));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4723_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12872 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_5 ), 
            .I2(\REG.mem_11_5 ), .I3(rd_addr_r[1]), .O(n15073));
    defparam rd_addr_r_0__bdd_4_lut_12872.LUT_INIT = 16'he4aa;
    SB_LUT4 i4219_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_2_31 ), .O(n5693));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4219_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4218_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_2_30 ), .O(n5692));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4218_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11117_3_lut (.I0(\REG.mem_20_14 ), .I1(\REG.mem_21_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13228));
    defparam i11117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11118_3_lut (.I0(\REG.mem_22_14 ), .I1(\REG.mem_23_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13229));
    defparam i11118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11115_3_lut (.I0(\REG.mem_18_14 ), .I1(\REG.mem_19_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13226));
    defparam i11115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11114_3_lut (.I0(\REG.mem_16_14 ), .I1(\REG.mem_17_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13225));
    defparam i11114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11522_3_lut (.I0(\REG.mem_20_26 ), .I1(\REG.mem_21_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13633));
    defparam i11522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11523_3_lut (.I0(\REG.mem_22_26 ), .I1(\REG.mem_23_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13634));
    defparam i11523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11105_3_lut (.I0(\REG.mem_4_14 ), .I1(\REG.mem_5_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13216));
    defparam i11105_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11106_3_lut (.I0(\REG.mem_6_14 ), .I1(\REG.mem_7_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13217));
    defparam i11106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11601_3_lut (.I0(\REG.mem_18_26 ), .I1(\REG.mem_19_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13712));
    defparam i11601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11600_3_lut (.I0(\REG.mem_16_26 ), .I1(\REG.mem_17_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13711));
    defparam i11600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11103_3_lut (.I0(\REG.mem_2_14 ), .I1(\REG.mem_3_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13214));
    defparam i11103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11102_3_lut (.I0(\REG.mem_0_14 ), .I1(\REG.mem_1_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13213));
    defparam i11102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11099_3_lut (.I0(n14584), .I1(n14524), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13210));
    defparam i11099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11435_3_lut (.I0(\REG.mem_20_3 ), .I1(\REG.mem_21_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13546));
    defparam i11435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11436_3_lut (.I0(\REG.mem_22_3 ), .I1(\REG.mem_23_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13547));
    defparam i11436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11636_3_lut (.I0(\REG.mem_12_27 ), .I1(\REG.mem_13_27 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13747));
    defparam i11636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11637_3_lut (.I0(\REG.mem_14_27 ), .I1(\REG.mem_15_27 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13748));
    defparam i11637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12024_3_lut (.I0(\REG.mem_10_27 ), .I1(\REG.mem_11_27 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14135));
    defparam i12024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12023_3_lut (.I0(\REG.mem_8_27 ), .I1(\REG.mem_9_27 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14134));
    defparam i12023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12051_3_lut (.I0(\REG.mem_18_3 ), .I1(\REG.mem_19_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14162));
    defparam i12051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12050_3_lut (.I0(\REG.mem_16_3 ), .I1(\REG.mem_17_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14161));
    defparam i12050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11225_3_lut (.I0(\REG.mem_4_29 ), .I1(\REG.mem_5_29 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13336));
    defparam i11225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11226_3_lut (.I0(\REG.mem_6_29 ), .I1(\REG.mem_7_29 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13337));
    defparam i11226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11733_3_lut (.I0(\REG.mem_2_29 ), .I1(\REG.mem_3_29 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13844));
    defparam i11733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11732_3_lut (.I0(\REG.mem_0_29 ), .I1(\REG.mem_1_29 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13843));
    defparam i11732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10997_3_lut (.I0(\REG.mem_20_30 ), .I1(\REG.mem_21_30 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13108));
    defparam i10997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10998_3_lut (.I0(\REG.mem_22_30 ), .I1(\REG.mem_23_30 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13109));
    defparam i10998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10986_3_lut (.I0(\REG.mem_18_30 ), .I1(\REG.mem_19_30 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13097));
    defparam i10986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10985_3_lut (.I0(\REG.mem_16_30 ), .I1(\REG.mem_17_30 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13096));
    defparam i10985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8021256_i1_3_lut (.I0(n14686), .I1(n16102), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[5]));
    defparam i8021256_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7823157_i1_3_lut (.I0(n15064), .I1(n15028), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[6]));
    defparam i7823157_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8621556_i1_3_lut (.I0(n13608), .I1(n14710), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[8]));
    defparam i8621556_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11497_3_lut (.I0(n15364), .I1(n13607), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n13608));
    defparam i11497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11496_3_lut (.I0(n15658), .I1(n15466), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13607));
    defparam i11496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7979235_i1_3_lut (.I0(n15340), .I1(n15304), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[13]));
    defparam i7979235_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8573532_i1_3_lut (.I0(n14530), .I1(n16222), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[16]));
    defparam i8573532_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8477484_i1_3_lut (.I0(n14656), .I1(n14974), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[19]));
    defparam i8477484_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8453472_i1_3_lut (.I0(n13560), .I1(n14560), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[20]));
    defparam i8453472_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11449_3_lut (.I0(n15166), .I1(n13559), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n13560));
    defparam i11449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11448_3_lut (.I0(n16018), .I1(n16000), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13559));
    defparam i11448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8429460_i1_3_lut (.I0(n16030), .I1(n16156), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[21]));
    defparam i8429460_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8357424_i1_3_lut (.I0(n15040), .I1(n14920), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[24]));
    defparam i8357424_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8333412_i1_3_lut (.I0(n15610), .I1(n15526), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[25]));
    defparam i8333412_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8261376_i1_3_lut (.I0(n13776), .I1(n14698), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[28]));
    defparam i8261376_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11665_3_lut (.I0(n15628), .I1(n13775), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n13776));
    defparam i11665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11664_3_lut (.I0(n15676), .I1(n15604), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13775));
    defparam i11664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wp_sync2_r_5__I_0_130_i1_2_lut (.I0(wp_sync2_r[4]), .I1(wp_sync2_r[5]), 
            .I2(GND_net), .I3(GND_net), .O(wp_sync_w[4]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam wp_sync2_r_5__I_0_130_i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i5_1_lut (.I0(rd_addr_r[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i4_1_lut (.I0(rd_addr_r[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i3_1_lut (.I0(rd_addr_r[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i2_1_lut (.I0(rd_addr_r[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i1_1_lut (.I0(rd_addr_r[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11624_3_lut (.I0(\REG.mem_4_15 ), .I1(\REG.mem_5_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13735));
    defparam i11624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11625_3_lut (.I0(\REG.mem_6_15 ), .I1(\REG.mem_7_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13736));
    defparam i11625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12069_3_lut (.I0(\REG.mem_2_15 ), .I1(\REG.mem_3_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14180));
    defparam i12069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12068_3_lut (.I0(\REG.mem_0_15 ), .I1(\REG.mem_1_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14179));
    defparam i12068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4217_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_2_29 ), .O(n5691));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4217_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut (.I0(wp_sync2_r[1]), .I1(wp_sync2_r[2]), .I2(wp_sync_w[3]), 
            .I3(GND_net), .O(wp_sync_w[1]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i12026_3_lut (.I0(\REG.mem_4_3 ), .I1(\REG.mem_5_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14137));
    defparam i12026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12027_3_lut (.I0(\REG.mem_6_3 ), .I1(\REG.mem_7_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14138));
    defparam i12027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12044_3_lut (.I0(\REG.mem_12_3 ), .I1(\REG.mem_13_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14155));
    defparam i12044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12045_3_lut (.I0(\REG.mem_14_3 ), .I1(\REG.mem_15_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14156));
    defparam i12045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12021_3_lut (.I0(\REG.mem_2_3 ), .I1(\REG.mem_3_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14132));
    defparam i12021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12020_3_lut (.I0(\REG.mem_0_3 ), .I1(\REG.mem_1_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14131));
    defparam i12020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_74 (.I0(wp_sync2_r[3]), .I1(wp_sync2_r[5]), 
            .I2(wp_sync2_r[4]), .I3(GND_net), .O(wp_sync_w[3]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_adj_74.LUT_INIT = 16'h9696;
    SB_LUT4 i12033_3_lut (.I0(\REG.mem_10_3 ), .I1(\REG.mem_11_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14144));
    defparam i12033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12032_3_lut (.I0(\REG.mem_8_3 ), .I1(\REG.mem_9_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14143));
    defparam i12032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4216_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_2_28 ), .O(n5690));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4216_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4215_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_2_27 ), .O(n5689));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4215_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4511_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_12_3 ), .O(n5985));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4511_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4510_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_12_2 ), .O(n5984));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4510_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4509_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_12_1 ), .O(n5983));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4509_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4508_3_lut_4_lut (.I0(n28_adj_1375), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_12_0 ), .O(n5982));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4508_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11010_3_lut (.I0(n14782), .I1(n15772), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13121));
    defparam i11010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_nxt_c_5__I_0_138_i4_2_lut (.I0(\rd_addr_nxt_c_5__N_573[3] ), 
            .I1(\rd_addr_nxt_c_5__N_573[4] ), .I2(GND_net), .I3(GND_net), 
            .O(rd_grey_w[3]));   // src/fifo_dc_32_lut_gen.v(504[28:66])
    defparam rd_addr_nxt_c_5__I_0_138_i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10988_3_lut (.I0(\REG.mem_20_11 ), .I1(\REG.mem_21_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13099));
    defparam i10988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10989_3_lut (.I0(\REG.mem_22_11 ), .I1(\REG.mem_23_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13100));
    defparam i10989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10980_3_lut (.I0(\REG.mem_18_11 ), .I1(\REG.mem_19_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13091));
    defparam i10980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10979_3_lut (.I0(\REG.mem_16_11 ), .I1(\REG.mem_17_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13090));
    defparam i10979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12005_3_lut (.I0(\REG.mem_28_4 ), .I1(\REG.mem_29_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14116));
    defparam i12005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12006_3_lut (.I0(\REG.mem_30_4 ), .I1(\REG.mem_31_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14117));
    defparam i12006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12000_3_lut (.I0(\REG.mem_26_4 ), .I1(\REG.mem_27_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14111));
    defparam i12000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11999_3_lut (.I0(\REG.mem_24_4 ), .I1(\REG.mem_25_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14110));
    defparam i11999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4214_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_2_26 ), .O(n5688));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4214_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4213_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_2_25 ), .O(n5687));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4213_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4212_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_2_24 ), .O(n5686));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4212_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4211_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_2_23 ), .O(n5685));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4211_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10958_3_lut (.I0(\REG.mem_4_11 ), .I1(\REG.mem_5_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13069));
    defparam i10958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10959_3_lut (.I0(\REG.mem_6_11 ), .I1(\REG.mem_7_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13070));
    defparam i10959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11300_3_lut (.I0(\REG.mem_28_1 ), .I1(\REG.mem_29_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13411));
    defparam i11300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11301_3_lut (.I0(\REG.mem_30_1 ), .I1(\REG.mem_31_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13412));
    defparam i11301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4210_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_2_22 ), .O(n5684));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4210_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4209_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_2_21 ), .O(n5683));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4209_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4208_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_2_20 ), .O(n5682));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4208_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4207_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_2_19 ), .O(n5681));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4207_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4206_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_2_18 ), .O(n5680));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4206_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4205_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_2_17 ), .O(n5679));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4205_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4204_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_2_16 ), .O(n5678));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4204_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11295_3_lut (.I0(\REG.mem_26_1 ), .I1(\REG.mem_27_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13406));
    defparam i11295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11294_3_lut (.I0(\REG.mem_24_1 ), .I1(\REG.mem_25_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13405));
    defparam i11294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4203_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_2_15 ), .O(n5677));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4203_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11498_3_lut (.I0(n14614), .I1(n14494), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13609));
    defparam i11498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11493_3_lut (.I0(n15238), .I1(n15184), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13604));
    defparam i11493_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4202_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_2_14 ), .O(n5676));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4202_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4201_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_2_13 ), .O(n5675));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4201_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4200_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_2_12 ), .O(n5674));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4200_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4087_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_0_6 ), .O(n5561));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4087_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_75 (.I0(rp_sync2_r[2]), .I1(rp_sync_w[3]), 
            .I2(rp_sync2_r[1]), .I3(GND_net), .O(rp_sync_w[1]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_3_lut_adj_75.LUT_INIT = 16'h9696;
    SB_LUT4 i4199_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_2_11 ), .O(n5673));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4199_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4198_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_2_10 ), .O(n5672));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4198_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11441_3_lut (.I0(\REG.mem_12_31 ), .I1(\REG.mem_13_31 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13552));
    defparam i11441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11442_3_lut (.I0(\REG.mem_14_31 ), .I1(\REG.mem_15_31 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13553));
    defparam i11442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11433_3_lut (.I0(\REG.mem_10_31 ), .I1(\REG.mem_11_31 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13544));
    defparam i11433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11432_3_lut (.I0(\REG.mem_8_31 ), .I1(\REG.mem_9_31 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13543));
    defparam i11432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11543_3_lut (.I0(\REG.mem_4_8 ), .I1(\REG.mem_5_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13654));
    defparam i11543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11544_3_lut (.I0(\REG.mem_6_8 ), .I1(\REG.mem_7_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13655));
    defparam i11544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11688_3_lut (.I0(\REG.mem_2_8 ), .I1(\REG.mem_3_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13799));
    defparam i11688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11687_3_lut (.I0(\REG.mem_0_8 ), .I1(\REG.mem_1_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13798));
    defparam i11687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12014_3_lut (.I0(\REG.mem_28_23 ), .I1(\REG.mem_29_23 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14125));
    defparam i12014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12015_3_lut (.I0(\REG.mem_30_23 ), .I1(\REG.mem_31_23 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14126));
    defparam i12015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12009_3_lut (.I0(\REG.mem_26_23 ), .I1(\REG.mem_27_23 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14120));
    defparam i12009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12008_3_lut (.I0(\REG.mem_24_23 ), .I1(\REG.mem_25_23 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14119));
    defparam i12008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11606_3_lut (.I0(\REG.mem_4_12 ), .I1(\REG.mem_5_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13717));
    defparam i11606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11607_3_lut (.I0(\REG.mem_6_12 ), .I1(\REG.mem_7_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13718));
    defparam i11607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11328_3_lut (.I0(\REG.mem_2_12 ), .I1(\REG.mem_3_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13439));
    defparam i11328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11327_3_lut (.I0(\REG.mem_0_12 ), .I1(\REG.mem_1_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13438));
    defparam i11327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11084_3_lut (.I0(\REG.mem_12_18 ), .I1(\REG.mem_13_18 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13195));
    defparam i11084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11085_3_lut (.I0(\REG.mem_14_18 ), .I1(\REG.mem_15_18 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13196));
    defparam i11085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11082_3_lut (.I0(\REG.mem_10_18 ), .I1(\REG.mem_11_18 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13193));
    defparam i11082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11081_3_lut (.I0(\REG.mem_8_18 ), .I1(\REG.mem_9_18 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13192));
    defparam i11081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11465_3_lut (.I0(\REG.mem_28_12 ), .I1(\REG.mem_29_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13576));
    defparam i11465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11466_3_lut (.I0(\REG.mem_30_12 ), .I1(\REG.mem_31_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13577));
    defparam i11466_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11439_3_lut (.I0(\REG.mem_26_12 ), .I1(\REG.mem_27_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13550));
    defparam i11439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11438_3_lut (.I0(\REG.mem_24_12 ), .I1(\REG.mem_25_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13549));
    defparam i11438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11024_3_lut (.I0(\REG.mem_28_17 ), .I1(\REG.mem_29_17 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13135));
    defparam i11024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11025_3_lut (.I0(\REG.mem_30_17 ), .I1(\REG.mem_31_17 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13136));
    defparam i11025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11016_3_lut (.I0(\REG.mem_26_17 ), .I1(\REG.mem_27_17 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13127));
    defparam i11016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11015_3_lut (.I0(\REG.mem_24_17 ), .I1(\REG.mem_25_17 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13126));
    defparam i11015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10943_3_lut (.I0(n16198), .I1(n16192), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13054));
    defparam i10943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10944_3_lut (.I0(n16174), .I1(n16150), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13055));
    defparam i10944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11471_3_lut (.I0(n14518), .I1(n16210), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13582));
    defparam i11471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11096_3_lut (.I0(\REG.mem_28_18 ), .I1(\REG.mem_29_18 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13207));
    defparam i11096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11097_3_lut (.I0(\REG.mem_30_18 ), .I1(\REG.mem_31_18 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13208));
    defparam i11097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11094_3_lut (.I0(\REG.mem_26_18 ), .I1(\REG.mem_27_18 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13205));
    defparam i11094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11093_3_lut (.I0(\REG.mem_24_18 ), .I1(\REG.mem_25_18 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13204));
    defparam i11093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11111_3_lut (.I0(\REG.mem_12_14 ), .I1(\REG.mem_13_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13222));
    defparam i11111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11112_3_lut (.I0(\REG.mem_14_14 ), .I1(\REG.mem_15_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13223));
    defparam i11112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4197_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_2_9 ), .O(n5671));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4197_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4196_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_2_8 ), .O(n5670));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4196_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4195_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_2_7 ), .O(n5669));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4195_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4194_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_2_6 ), .O(n5668));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4194_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4193_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_2_5 ), .O(n5667));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4193_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11109_3_lut (.I0(\REG.mem_10_14 ), .I1(\REG.mem_11_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13220));
    defparam i11109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11108_3_lut (.I0(\REG.mem_8_14 ), .I1(\REG.mem_9_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13219));
    defparam i11108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11123_3_lut (.I0(\REG.mem_28_14 ), .I1(\REG.mem_29_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13234));
    defparam i11123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11124_3_lut (.I0(\REG.mem_30_14 ), .I1(\REG.mem_31_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13235));
    defparam i11124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11121_3_lut (.I0(\REG.mem_26_14 ), .I1(\REG.mem_27_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13232));
    defparam i11121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11120_3_lut (.I0(\REG.mem_24_14 ), .I1(\REG.mem_25_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13231));
    defparam i11120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11483_3_lut (.I0(\REG.mem_12_26 ), .I1(\REG.mem_13_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13594));
    defparam i11483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11484_3_lut (.I0(\REG.mem_14_26 ), .I1(\REG.mem_15_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13595));
    defparam i11484_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11451_3_lut (.I0(\REG.mem_10_26 ), .I1(\REG.mem_11_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13562));
    defparam i11451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11450_3_lut (.I0(\REG.mem_8_26 ), .I1(\REG.mem_9_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13561));
    defparam i11450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11144_3_lut (.I0(\REG.mem_12_9 ), .I1(\REG.mem_13_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13255));
    defparam i11144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11145_3_lut (.I0(\REG.mem_14_9 ), .I1(\REG.mem_15_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13256));
    defparam i11145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11139_3_lut (.I0(\REG.mem_10_9 ), .I1(\REG.mem_11_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13250));
    defparam i11139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11138_3_lut (.I0(\REG.mem_8_9 ), .I1(\REG.mem_9_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13249));
    defparam i11138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12104_3_lut (.I0(\REG.mem_4_20 ), .I1(\REG.mem_5_20 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14215));
    defparam i12104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12105_3_lut (.I0(\REG.mem_6_20 ), .I1(\REG.mem_7_20 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14216));
    defparam i12105_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12102_3_lut (.I0(\REG.mem_2_20 ), .I1(\REG.mem_3_20 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14213));
    defparam i12102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12101_3_lut (.I0(\REG.mem_0_20 ), .I1(\REG.mem_1_20 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14212));
    defparam i12101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12047_3_lut (.I0(n14536), .I1(n16216), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n14158));
    defparam i12047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12030_3_lut (.I0(n14644), .I1(n14596), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n14141));
    defparam i12030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12029_3_lut (.I0(n14728), .I1(n14668), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n14140));
    defparam i12029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11585_3_lut (.I0(\REG.mem_28_26 ), .I1(\REG.mem_29_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13696));
    defparam i11585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11586_3_lut (.I0(\REG.mem_30_26 ), .I1(\REG.mem_31_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13697));
    defparam i11586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11532_3_lut (.I0(\REG.mem_26_26 ), .I1(\REG.mem_27_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13643));
    defparam i11532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11531_3_lut (.I0(\REG.mem_24_26 ), .I1(\REG.mem_25_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13642));
    defparam i11531_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11456_3_lut (.I0(n14500), .I1(n16228), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n13567));
    defparam i11456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12018_3_lut (.I0(n14578), .I1(n14554), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n14129));
    defparam i12018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12017_3_lut (.I0(n16114), .I1(n14620), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n14128));
    defparam i12017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11150_3_lut (.I0(\REG.mem_12_7 ), .I1(\REG.mem_13_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13261));
    defparam i11150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11151_3_lut (.I0(\REG.mem_14_7 ), .I1(\REG.mem_15_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13262));
    defparam i11151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11142_3_lut (.I0(\REG.mem_10_7 ), .I1(\REG.mem_11_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13253));
    defparam i11142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11141_3_lut (.I0(\REG.mem_8_7 ), .I1(\REG.mem_9_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13252));
    defparam i11141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4192_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_2_4 ), .O(n5666));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4192_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11090_3_lut (.I0(\REG.mem_20_18 ), .I1(\REG.mem_21_18 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13201));
    defparam i11090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11091_3_lut (.I0(\REG.mem_22_18 ), .I1(\REG.mem_23_18 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13202));
    defparam i11091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11088_3_lut (.I0(\REG.mem_18_18 ), .I1(\REG.mem_19_18 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13199));
    defparam i11088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11087_3_lut (.I0(\REG.mem_16_18 ), .I1(\REG.mem_17_18 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13198));
    defparam i11087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11000_3_lut (.I0(\REG.mem_28_11 ), .I1(\REG.mem_29_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13111));
    defparam i11000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11001_3_lut (.I0(\REG.mem_30_11 ), .I1(\REG.mem_31_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13112));
    defparam i11001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10995_3_lut (.I0(\REG.mem_26_11 ), .I1(\REG.mem_27_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13106));
    defparam i10995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10994_3_lut (.I0(\REG.mem_24_11 ), .I1(\REG.mem_25_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13105));
    defparam i10994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4153_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_2_1 ), .O(n5627));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4153_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11513_3_lut (.I0(\REG.mem_28_29 ), .I1(\REG.mem_29_29 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13624));
    defparam i11513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11514_3_lut (.I0(\REG.mem_30_29 ), .I1(\REG.mem_31_29 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13625));
    defparam i11514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11481_3_lut (.I0(\REG.mem_26_29 ), .I1(\REG.mem_27_29 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13592));
    defparam i11481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11480_3_lut (.I0(\REG.mem_24_29 ), .I1(\REG.mem_25_29 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13591));
    defparam i11480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11174_3_lut (.I0(\REG.mem_28_7 ), .I1(\REG.mem_29_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13285));
    defparam i11174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11175_3_lut (.I0(\REG.mem_30_7 ), .I1(\REG.mem_31_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13286));
    defparam i11175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11172_3_lut (.I0(\REG.mem_26_7 ), .I1(\REG.mem_27_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13283));
    defparam i11172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11171_3_lut (.I0(\REG.mem_24_7 ), .I1(\REG.mem_25_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13282));
    defparam i11171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11546_3_lut (.I0(\REG.mem_28_15 ), .I1(\REG.mem_29_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13657));
    defparam i11546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11547_3_lut (.I0(\REG.mem_30_15 ), .I1(\REG.mem_31_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13658));
    defparam i11547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4152_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_2_0 ), .O(n5626));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4152_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4166_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_2_2 ), .O(n5640));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4166_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4176_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_2_3 ), .O(n5650));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4176_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11505_3_lut (.I0(\REG.mem_26_15 ), .I1(\REG.mem_27_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13616));
    defparam i11505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11504_3_lut (.I0(\REG.mem_24_15 ), .I1(\REG.mem_25_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13615));
    defparam i11504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i10_2_lut_3_lut_4_lut (.I0(dc32_fifo_write_enable), 
            .I1(dc32_fifo_full), .I2(\wr_addr_r[0] ), .I3(wr_addr_r[1]), 
            .O(n10_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i10_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i11189_3_lut (.I0(\REG.mem_12_10 ), .I1(\REG.mem_13_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13300));
    defparam i11189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11190_3_lut (.I0(\REG.mem_14_10 ), .I1(\REG.mem_15_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13301));
    defparam i11190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i8_2_lut_3_lut_4_lut (.I0(dc32_fifo_write_enable), 
            .I1(dc32_fifo_full), .I2(\wr_addr_r[0] ), .I3(wr_addr_r[1]), 
            .O(n8_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i8_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i11187_3_lut (.I0(\REG.mem_10_10 ), .I1(\REG.mem_11_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13298));
    defparam i11187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11186_3_lut (.I0(\REG.mem_8_10 ), .I1(\REG.mem_9_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13297));
    defparam i11186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11153_3_lut (.I0(\REG.mem_20_9 ), .I1(\REG.mem_21_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13264));
    defparam i11153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11154_3_lut (.I0(\REG.mem_22_9 ), .I1(\REG.mem_23_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13265));
    defparam i11154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11148_3_lut (.I0(\REG.mem_18_9 ), .I1(\REG.mem_19_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13259));
    defparam i11148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11147_3_lut (.I0(\REG.mem_16_9 ), .I1(\REG.mem_17_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13258));
    defparam i11147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11264_3_lut (.I0(\REG.mem_28_2 ), .I1(\REG.mem_29_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13375));
    defparam i11264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11265_3_lut (.I0(\REG.mem_30_2 ), .I1(\REG.mem_31_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13376));
    defparam i11265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11259_3_lut (.I0(\REG.mem_26_2 ), .I1(\REG.mem_27_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13370));
    defparam i11259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11258_3_lut (.I0(\REG.mem_24_2 ), .I1(\REG.mem_25_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13369));
    defparam i11258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11750_3_lut (.I0(\REG.mem_28_30 ), .I1(\REG.mem_29_30 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13861));
    defparam i11750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11751_3_lut (.I0(\REG.mem_30_30 ), .I1(\REG.mem_31_30 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13862));
    defparam i11751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11007_3_lut (.I0(\REG.mem_26_30 ), .I1(\REG.mem_27_30 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13118));
    defparam i11007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11006_3_lut (.I0(\REG.mem_24_30 ), .I1(\REG.mem_25_30 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n13117));
    defparam i11006_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module FIFO_Quad_Word
//

module FIFO_Quad_Word (n8, rd_addr_r, SLM_CLK_c, reset_all_w, wr_addr_r, 
            rx_buf_byte, n4446, GND_net, \wr_addr_p1_w[2] , n12215, 
            rd_fifo_en_w, \mem_LUT.data_raw_r[0] , n8_adj_2, n5599, 
            n5607, n12439, VCC_net, is_tx_fifo_full_flag, n5645, \fifo_temp_output[7] , 
            n5648, \fifo_temp_output[6] , n5653, \fifo_temp_output[5] , 
            n6947, \fifo_temp_output[0] , n5656, \fifo_temp_output[4] , 
            n5659, \fifo_temp_output[3] , n5662, \fifo_temp_output[2] , 
            n5665, \fifo_temp_output[1] , n6923, n6920, fifo_write_cmd, 
            wr_fifo_en_w, n5636, rd_fifo_en_prev_r, \mem_LUT.data_raw_r[1] , 
            \mem_LUT.data_raw_r[2] , \mem_LUT.data_raw_r[3] , \mem_LUT.data_raw_r[4] , 
            \mem_LUT.data_raw_r[5] , \mem_LUT.data_raw_r[6] , \mem_LUT.data_raw_r[7] , 
            n12836, is_fifo_empty_flag, fifo_read_cmd, \rd_addr_p1_w[2] , 
            \rd_addr_p1_w[1] ) /* synthesis syn_module_defined=1 */ ;
    input n8;
    output [2:0]rd_addr_r;
    input SLM_CLK_c;
    input reset_all_w;
    output [2:0]wr_addr_r;
    input [7:0]rx_buf_byte;
    output n4446;
    input GND_net;
    output \wr_addr_p1_w[2] ;
    output n12215;
    output rd_fifo_en_w;
    output \mem_LUT.data_raw_r[0] ;
    input n8_adj_2;
    input n5599;
    input n5607;
    input n12439;
    input VCC_net;
    output is_tx_fifo_full_flag;
    input n5645;
    output \fifo_temp_output[7] ;
    input n5648;
    output \fifo_temp_output[6] ;
    input n5653;
    output \fifo_temp_output[5] ;
    input n6947;
    output \fifo_temp_output[0] ;
    input n5656;
    output \fifo_temp_output[4] ;
    input n5659;
    output \fifo_temp_output[3] ;
    input n5662;
    output \fifo_temp_output[2] ;
    input n5665;
    output \fifo_temp_output[1] ;
    input n6923;
    input n6920;
    input fifo_write_cmd;
    output wr_fifo_en_w;
    input n5636;
    output rd_fifo_en_prev_r;
    output \mem_LUT.data_raw_r[1] ;
    output \mem_LUT.data_raw_r[2] ;
    output \mem_LUT.data_raw_r[3] ;
    output \mem_LUT.data_raw_r[4] ;
    output \mem_LUT.data_raw_r[5] ;
    output \mem_LUT.data_raw_r[6] ;
    output \mem_LUT.data_raw_r[7] ;
    input n12836;
    output is_fifo_empty_flag;
    input fifo_read_cmd;
    output \rd_addr_p1_w[2] ;
    output \rd_addr_p1_w[1] ;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_3 lscc_fifo_inst (.n8(n8), 
            .rd_addr_r({rd_addr_r}), .SLM_CLK_c(SLM_CLK_c), .reset_all_w(reset_all_w), 
            .wr_addr_r({wr_addr_r}), .rx_buf_byte({rx_buf_byte}), .n4446(n4446), 
            .GND_net(GND_net), .\wr_addr_p1_w[2] (\wr_addr_p1_w[2] ), .n12215(n12215), 
            .rd_fifo_en_w(rd_fifo_en_w), .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r[0] ), 
            .n8_adj_1(n8_adj_2), .n5599(n5599), .n5607(n5607), .n12439(n12439), 
            .VCC_net(VCC_net), .is_tx_fifo_full_flag(is_tx_fifo_full_flag), 
            .n5645(n5645), .\fifo_temp_output[7] (\fifo_temp_output[7] ), 
            .n5648(n5648), .\fifo_temp_output[6] (\fifo_temp_output[6] ), 
            .n5653(n5653), .\fifo_temp_output[5] (\fifo_temp_output[5] ), 
            .n6947(n6947), .\fifo_temp_output[0] (\fifo_temp_output[0] ), 
            .n5656(n5656), .\fifo_temp_output[4] (\fifo_temp_output[4] ), 
            .n5659(n5659), .\fifo_temp_output[3] (\fifo_temp_output[3] ), 
            .n5662(n5662), .\fifo_temp_output[2] (\fifo_temp_output[2] ), 
            .n5665(n5665), .\fifo_temp_output[1] (\fifo_temp_output[1] ), 
            .n6923(n6923), .n6920(n6920), .fifo_write_cmd(fifo_write_cmd), 
            .wr_fifo_en_w(wr_fifo_en_w), .n5636(n5636), .rd_fifo_en_prev_r(rd_fifo_en_prev_r), 
            .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r[1] ), .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r[2] ), 
            .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r[3] ), .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r[4] ), 
            .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r[5] ), .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r[6] ), 
            .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r[7] ), .n12836(n12836), 
            .is_fifo_empty_flag(is_fifo_empty_flag), .fifo_read_cmd(fifo_read_cmd), 
            .\rd_addr_p1_w[2] (\rd_addr_p1_w[2] ), .\rd_addr_p1_w[1] (\rd_addr_p1_w[1] )) /* synthesis syn_module_defined=1 */ ;   // src/fifo_quad_word_mod.v(20[37:380])
    
endmodule
//
// Verilog Description of module FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_3
//

module FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_3 (n8, 
            rd_addr_r, SLM_CLK_c, reset_all_w, wr_addr_r, rx_buf_byte, 
            n4446, GND_net, \wr_addr_p1_w[2] , n12215, rd_fifo_en_w, 
            \mem_LUT.data_raw_r[0] , n8_adj_1, n5599, n5607, n12439, 
            VCC_net, is_tx_fifo_full_flag, n5645, \fifo_temp_output[7] , 
            n5648, \fifo_temp_output[6] , n5653, \fifo_temp_output[5] , 
            n6947, \fifo_temp_output[0] , n5656, \fifo_temp_output[4] , 
            n5659, \fifo_temp_output[3] , n5662, \fifo_temp_output[2] , 
            n5665, \fifo_temp_output[1] , n6923, n6920, fifo_write_cmd, 
            wr_fifo_en_w, n5636, rd_fifo_en_prev_r, \mem_LUT.data_raw_r[1] , 
            \mem_LUT.data_raw_r[2] , \mem_LUT.data_raw_r[3] , \mem_LUT.data_raw_r[4] , 
            \mem_LUT.data_raw_r[5] , \mem_LUT.data_raw_r[6] , \mem_LUT.data_raw_r[7] , 
            n12836, is_fifo_empty_flag, fifo_read_cmd, \rd_addr_p1_w[2] , 
            \rd_addr_p1_w[1] ) /* synthesis syn_module_defined=1 */ ;
    input n8;
    output [2:0]rd_addr_r;
    input SLM_CLK_c;
    input reset_all_w;
    output [2:0]wr_addr_r;
    input [7:0]rx_buf_byte;
    output n4446;
    input GND_net;
    output \wr_addr_p1_w[2] ;
    output n12215;
    output rd_fifo_en_w;
    output \mem_LUT.data_raw_r[0] ;
    input n8_adj_1;
    input n5599;
    input n5607;
    input n12439;
    input VCC_net;
    output is_tx_fifo_full_flag;
    input n5645;
    output \fifo_temp_output[7] ;
    input n5648;
    output \fifo_temp_output[6] ;
    input n5653;
    output \fifo_temp_output[5] ;
    input n6947;
    output \fifo_temp_output[0] ;
    input n5656;
    output \fifo_temp_output[4] ;
    input n5659;
    output \fifo_temp_output[3] ;
    input n5662;
    output \fifo_temp_output[2] ;
    input n5665;
    output \fifo_temp_output[1] ;
    input n6923;
    input n6920;
    input fifo_write_cmd;
    output wr_fifo_en_w;
    input n5636;
    output rd_fifo_en_prev_r;
    output \mem_LUT.data_raw_r[1] ;
    output \mem_LUT.data_raw_r[2] ;
    output \mem_LUT.data_raw_r[3] ;
    output \mem_LUT.data_raw_r[4] ;
    output \mem_LUT.data_raw_r[5] ;
    output \mem_LUT.data_raw_r[6] ;
    output \mem_LUT.data_raw_r[7] ;
    input n12836;
    output is_fifo_empty_flag;
    input fifo_read_cmd;
    output \rd_addr_p1_w[2] ;
    output \rd_addr_p1_w[1] ;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n3, \mem_LUT.mem_3_7 , n6917, n2, \mem_LUT.mem_3_6 , n6916, 
        \mem_LUT.mem_3_5 , n6915, \mem_LUT.mem_3_4 , n6914, \mem_LUT.mem_3_3 , 
        n6913, \mem_LUT.mem_3_2 , n6912, \mem_LUT.mem_3_1 , n6911, 
        \mem_LUT.mem_3_0 , n6910, n4, \mem_LUT.mem_2_7 , n6901, \mem_LUT.mem_2_6 , 
        n6900, \mem_LUT.mem_2_5 , n6899, \mem_LUT.mem_2_4 , n6898, 
        \mem_LUT.mem_2_3 , n6897, \mem_LUT.mem_2_2 , n6896, \mem_LUT.mem_2_1 , 
        n6895, \mem_LUT.mem_2_0 , n6894, \mem_LUT.mem_1_7 , n6893, 
        \mem_LUT.mem_1_6 , n6892, \mem_LUT.mem_1_5 , n6891;
    wire [31:0]\mem_LUT.data_raw_r_31__N_1269 ;
    
    wire \mem_LUT.mem_1_4 , n6890, \mem_LUT.mem_1_3 , n6889, \mem_LUT.mem_1_2 , 
        n6888, \mem_LUT.mem_1_1 , n6887, \mem_LUT.mem_1_0 , n6886, 
        \mem_LUT.mem_0_7 , n6885, \mem_LUT.mem_0_6 , n6884, \mem_LUT.mem_0_5 , 
        n6883, \mem_LUT.mem_0_4 , n6882, \mem_LUT.mem_0_3 , n6881, 
        \mem_LUT.mem_0_2 , n6880, \mem_LUT.mem_0_1 , n6879, \mem_LUT.mem_0_0 , 
        n6878, n16165, n16123, n16117, n16093, n16081, n16069, 
        n16045, n16033;
    
    SB_DFFSR rd_addr_r__i0 (.Q(rd_addr_r[0]), .C(SLM_CLK_c), .D(n8), .R(reset_all_w));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 i5443_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_3_7 ), .O(n6917));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5443_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut (.I0(wr_addr_r[0]), .I1(rd_addr_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4446));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut (.I0(n4446), .I1(\wr_addr_p1_w[2] ), .I2(n2), .I3(rd_addr_r[2]), 
            .O(n12215));
    defparam i1_4_lut.LUT_INIT = 16'h0208;
    SB_LUT4 i5442_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_3_6 ), .O(n6916));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5442_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5441_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_3_5 ), .O(n6915));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5441_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5440_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_3_4 ), .O(n6914));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5440_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5439_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_3_3 ), .O(n6913));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5439_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5438_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_3_2 ), .O(n6912));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5438_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5437_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_3_1 ), .O(n6911));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5437_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5436_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_3_0 ), .O(n6910));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5436_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5427_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_2_7 ), .O(n6901));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5427_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5426_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_2_6 ), .O(n6900));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5426_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5425_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_2_5 ), .O(n6899));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5425_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5424_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_2_4 ), .O(n6898));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5424_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5423_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_2_3 ), .O(n6897));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5423_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5422_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_2_2 ), .O(n6896));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5422_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5421_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_2_1 ), .O(n6895));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5421_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5420_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_2_0 ), .O(n6894));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5420_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5419_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_1_7 ), .O(n6893));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5419_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5418_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_1_6 ), .O(n6892));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5418_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5417_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_1_5 ), .O(n6891));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5417_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \mem_LUT.data_raw_r__i1  (.Q(\mem_LUT.data_raw_r[0] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1269 [0]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_LUT4 i5416_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_1_4 ), .O(n6890));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5416_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5415_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_1_3 ), .O(n6889));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5415_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5414_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_1_2 ), .O(n6888));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5414_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5413_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_1_1 ), .O(n6887));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5413_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5412_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_1_0 ), .O(n6886));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5412_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5411_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_0_7 ), .O(n6885));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5411_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5410_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_0_6 ), .O(n6884));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5410_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5409_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_0_5 ), .O(n6883));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5409_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5408_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_0_4 ), .O(n6882));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5408_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5407_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_0_3 ), .O(n6881));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5407_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5406_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_0_2 ), .O(n6880));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5406_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5405_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_0_1 ), .O(n6879));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5405_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5404_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_0_0 ), .O(n6878));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5404_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFSR wr_addr_r__i0 (.Q(wr_addr_r[0]), .C(SLM_CLK_c), .D(n8_adj_1), 
            .R(reset_all_w));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 wr_addr_p1_w_1__I_0_i2_2_lut_3_lut (.I0(wr_addr_r[1]), .I1(wr_addr_r[0]), 
            .I2(rd_addr_r[1]), .I3(GND_net), .O(n2));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam wr_addr_p1_w_1__I_0_i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_DFF wr_addr_r__i2 (.Q(wr_addr_r[2]), .C(SLM_CLK_c), .D(n5599));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF wr_addr_r__i1 (.Q(wr_addr_r[1]), .C(SLM_CLK_c), .D(n5607));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFE full_r_84 (.Q(is_tx_fifo_full_flag), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n12439));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF \mem_LUT.data_buff_r__i7  (.Q(\fifo_temp_output[7] ), .C(SLM_CLK_c), 
           .D(n5645));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i6  (.Q(\fifo_temp_output[6] ), .C(SLM_CLK_c), 
           .D(n5648));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i5  (.Q(\fifo_temp_output[5] ), .C(SLM_CLK_c), 
           .D(n5653));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE \mem_LUT.data_buff_r__i0  (.Q(\fifo_temp_output[0] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n6947));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i4  (.Q(\fifo_temp_output[4] ), .C(SLM_CLK_c), 
           .D(n5656));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i3  (.Q(\fifo_temp_output[3] ), .C(SLM_CLK_c), 
           .D(n5659));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i2  (.Q(\fifo_temp_output[2] ), .C(SLM_CLK_c), 
           .D(n5662));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i1  (.Q(\fifo_temp_output[1] ), .C(SLM_CLK_c), 
           .D(n5665));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE rd_addr_r__i1 (.Q(rd_addr_r[1]), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n6923));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFE rd_addr_r__i2 (.Q(rd_addr_r[2]), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n6920));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF i347_348 (.Q(\mem_LUT.mem_3_7 ), .C(SLM_CLK_c), .D(n6917));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i344_345 (.Q(\mem_LUT.mem_3_6 ), .C(SLM_CLK_c), .D(n6916));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i341_342 (.Q(\mem_LUT.mem_3_5 ), .C(SLM_CLK_c), .D(n6915));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i338_339 (.Q(\mem_LUT.mem_3_4 ), .C(SLM_CLK_c), .D(n6914));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i335_336 (.Q(\mem_LUT.mem_3_3 ), .C(SLM_CLK_c), .D(n6913));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i332_333 (.Q(\mem_LUT.mem_3_2 ), .C(SLM_CLK_c), .D(n6912));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i329_330 (.Q(\mem_LUT.mem_3_1 ), .C(SLM_CLK_c), .D(n6911));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i326_327 (.Q(\mem_LUT.mem_3_0 ), .C(SLM_CLK_c), .D(n6910));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i251_252 (.Q(\mem_LUT.mem_2_7 ), .C(SLM_CLK_c), .D(n6901));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i248_249 (.Q(\mem_LUT.mem_2_6 ), .C(SLM_CLK_c), .D(n6900));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i245_246 (.Q(\mem_LUT.mem_2_5 ), .C(SLM_CLK_c), .D(n6899));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i242_243 (.Q(\mem_LUT.mem_2_4 ), .C(SLM_CLK_c), .D(n6898));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i239_240 (.Q(\mem_LUT.mem_2_3 ), .C(SLM_CLK_c), .D(n6897));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i236_237 (.Q(\mem_LUT.mem_2_2 ), .C(SLM_CLK_c), .D(n6896));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i233_234 (.Q(\mem_LUT.mem_2_1 ), .C(SLM_CLK_c), .D(n6895));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i230_231 (.Q(\mem_LUT.mem_2_0 ), .C(SLM_CLK_c), .D(n6894));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i155_156 (.Q(\mem_LUT.mem_1_7 ), .C(SLM_CLK_c), .D(n6893));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i152_153 (.Q(\mem_LUT.mem_1_6 ), .C(SLM_CLK_c), .D(n6892));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i149_150 (.Q(\mem_LUT.mem_1_5 ), .C(SLM_CLK_c), .D(n6891));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i146_147 (.Q(\mem_LUT.mem_1_4 ), .C(SLM_CLK_c), .D(n6890));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i143_144 (.Q(\mem_LUT.mem_1_3 ), .C(SLM_CLK_c), .D(n6889));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i140_141 (.Q(\mem_LUT.mem_1_2 ), .C(SLM_CLK_c), .D(n6888));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i137_138 (.Q(\mem_LUT.mem_1_1 ), .C(SLM_CLK_c), .D(n6887));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i134_135 (.Q(\mem_LUT.mem_1_0 ), .C(SLM_CLK_c), .D(n6886));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i59_60 (.Q(\mem_LUT.mem_0_7 ), .C(SLM_CLK_c), .D(n6885));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i56_57 (.Q(\mem_LUT.mem_0_6 ), .C(SLM_CLK_c), .D(n6884));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i53_54 (.Q(\mem_LUT.mem_0_5 ), .C(SLM_CLK_c), .D(n6883));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i50_51 (.Q(\mem_LUT.mem_0_4 ), .C(SLM_CLK_c), .D(n6882));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i47_48 (.Q(\mem_LUT.mem_0_3 ), .C(SLM_CLK_c), .D(n6881));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i44_45 (.Q(\mem_LUT.mem_0_2 ), .C(SLM_CLK_c), .D(n6880));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i41_42 (.Q(\mem_LUT.mem_0_1 ), .C(SLM_CLK_c), .D(n6879));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i38_39 (.Q(\mem_LUT.mem_0_0 ), .C(SLM_CLK_c), .D(n6878));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 i1709_3_lut (.I0(wr_addr_r[2]), .I1(wr_addr_r[1]), .I2(wr_addr_r[0]), 
            .I3(GND_net), .O(\wr_addr_p1_w[2] ));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam i1709_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 wr_en_i_I_0_2_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(GND_net), .I3(GND_net), .O(wr_fifo_en_w));   // src/fifo_quad_word_mod.v(103[21:60])
    defparam wr_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_DFF rd_fifo_en_prev_r_86 (.Q(rd_fifo_en_prev_r), .C(SLM_CLK_c), .D(n5636));   // src/fifo_quad_word_mod.v(353[29] 363[32])
    SB_DFFE \mem_LUT.data_raw_r__i2  (.Q(\mem_LUT.data_raw_r[1] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1269 [1]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i3  (.Q(\mem_LUT.data_raw_r[2] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1269 [2]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i4  (.Q(\mem_LUT.data_raw_r[3] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1269 [3]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i5  (.Q(\mem_LUT.data_raw_r[4] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1269 [4]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i6  (.Q(\mem_LUT.data_raw_r[5] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1269 [5]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i7  (.Q(\mem_LUT.data_raw_r[6] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1269 [6]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i8  (.Q(\mem_LUT.data_raw_r[7] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1269 [7]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_7 ), 
            .I2(\mem_LUT.mem_3_7 ), .I3(rd_addr_r[1]), .O(n16165));
    defparam rd_addr_r_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n16165_bdd_4_lut (.I0(n16165), .I1(\mem_LUT.mem_1_7 ), .I2(\mem_LUT.mem_0_7 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1269 [7]));
    defparam n16165_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13770 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_0 ), 
            .I2(\mem_LUT.mem_3_0 ), .I3(rd_addr_r[1]), .O(n16123));
    defparam rd_addr_r_0__bdd_4_lut_13770.LUT_INIT = 16'he4aa;
    SB_LUT4 n16123_bdd_4_lut (.I0(n16123), .I1(\mem_LUT.mem_1_0 ), .I2(\mem_LUT.mem_0_0 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1269 [0]));
    defparam n16123_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13735 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_6 ), 
            .I2(\mem_LUT.mem_3_6 ), .I3(rd_addr_r[1]), .O(n16117));
    defparam rd_addr_r_0__bdd_4_lut_13735.LUT_INIT = 16'he4aa;
    SB_LUT4 n16117_bdd_4_lut (.I0(n16117), .I1(\mem_LUT.mem_1_6 ), .I2(\mem_LUT.mem_0_6 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1269 [6]));
    defparam n16117_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13730 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_5 ), 
            .I2(\mem_LUT.mem_3_5 ), .I3(rd_addr_r[1]), .O(n16093));
    defparam rd_addr_r_0__bdd_4_lut_13730.LUT_INIT = 16'he4aa;
    SB_LUT4 n16093_bdd_4_lut (.I0(n16093), .I1(\mem_LUT.mem_1_5 ), .I2(\mem_LUT.mem_0_5 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1269 [5]));
    defparam n16093_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13710 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_4 ), 
            .I2(\mem_LUT.mem_3_4 ), .I3(rd_addr_r[1]), .O(n16081));
    defparam rd_addr_r_0__bdd_4_lut_13710.LUT_INIT = 16'he4aa;
    SB_LUT4 n16081_bdd_4_lut (.I0(n16081), .I1(\mem_LUT.mem_1_4 ), .I2(\mem_LUT.mem_0_4 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1269 [4]));
    defparam n16081_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13700 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_3 ), 
            .I2(\mem_LUT.mem_3_3 ), .I3(rd_addr_r[1]), .O(n16069));
    defparam rd_addr_r_0__bdd_4_lut_13700.LUT_INIT = 16'he4aa;
    SB_DFF empty_r_85 (.Q(is_fifo_empty_flag), .C(SLM_CLK_c), .D(n12836));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 n16069_bdd_4_lut (.I0(n16069), .I1(\mem_LUT.mem_1_3 ), .I2(\mem_LUT.mem_0_3 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1269 [3]));
    defparam n16069_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13690 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_2 ), 
            .I2(\mem_LUT.mem_3_2 ), .I3(rd_addr_r[1]), .O(n16045));
    defparam rd_addr_r_0__bdd_4_lut_13690.LUT_INIT = 16'he4aa;
    SB_LUT4 n16045_bdd_4_lut (.I0(n16045), .I1(\mem_LUT.mem_1_2 ), .I2(\mem_LUT.mem_0_2 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1269 [2]));
    defparam n16045_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_13670 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_1 ), 
            .I2(\mem_LUT.mem_3_1 ), .I3(rd_addr_r[1]), .O(n16033));
    defparam rd_addr_r_0__bdd_4_lut_13670.LUT_INIT = 16'he4aa;
    SB_LUT4 n16033_bdd_4_lut (.I0(n16033), .I1(\mem_LUT.mem_1_1 ), .I2(\mem_LUT.mem_0_1 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1269 [1]));
    defparam n16033_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_en_i_I_0_2_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(GND_net), .I3(GND_net), .O(rd_fifo_en_w));   // src/fifo_quad_word_mod.v(62[29:51])
    defparam rd_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1731_3_lut (.I0(rd_addr_r[2]), .I1(rd_addr_r[1]), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(\rd_addr_p1_w[2] ));   // src/fifo_quad_word_mod.v(71[47:65])
    defparam i1731_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1724_2_lut (.I0(rd_addr_r[1]), .I1(rd_addr_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(\rd_addr_p1_w[1] ));   // src/fifo_quad_word_mod.v(71[47:65])
    defparam i1724_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 EnabledDecoder_2_i3_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(GND_net), .O(n3));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i3_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i4_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(GND_net), .O(n4));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i4_2_lut_3_lut.LUT_INIT = 16'h0202;
>>>>>>> Stashed changes
>>>>>>> master
    
endmodule
//
// Verilog Description of module fifo_sc_32_lut_gen
//

<<<<<<< HEAD
module fifo_sc_32_lut_gen (SLM_CLK_c, sc32_fifo_almost_empty, reset_all, 
            GND_net, dc32_fifo_read_enable, sc32_fifo_read_enable) /* synthesis syn_module_defined=1 */ ;
    input SLM_CLK_c;
    output sc32_fifo_almost_empty;
    input reset_all;
    input GND_net;
    input dc32_fifo_read_enable;
    input sc32_fifo_read_enable;
=======
<<<<<<< Updated upstream
module clock (GND_net, VCC_net, ICE_SYSCLK_c, pll_clk_unbuf) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    input ICE_SYSCLK_c;
    output pll_clk_unbuf;
=======
module fifo_sc_32_lut_gen (DEBUG_9_c_0, SLM_CLK_c, \dc32_fifo_data_out[31] , 
            \dc32_fifo_data_out[30] , \dc32_fifo_data_out[29] , \dc32_fifo_data_out[28] , 
            \dc32_fifo_data_out[27] , \dc32_fifo_data_out[26] , \dc32_fifo_data_out[25] , 
            \dc32_fifo_data_out[24] , \dc32_fifo_data_out[23] , sc32_fifo_almost_empty, 
            reset_all, \dc32_fifo_data_out[22] , \dc32_fifo_data_out[21] , 
            \dc32_fifo_data_out[20] , \dc32_fifo_data_out[19] , \dc32_fifo_data_out[18] , 
            \dc32_fifo_data_out[17] , \dc32_fifo_data_out[16] , \dc32_fifo_data_out[15] , 
            \dc32_fifo_data_out[14] , \dc32_fifo_data_out[13] , \dc32_fifo_data_out[12] , 
            \dc32_fifo_data_out[11] , \dc32_fifo_data_out[10] , \dc32_fifo_data_out[9] , 
            \dc32_fifo_data_out[8] , \dc32_fifo_data_out[7] , \dc32_fifo_data_out[6] , 
            GND_net, \dc32_fifo_data_out[5] , \dc32_fifo_data_out[4] , 
            \dc32_fifo_data_out[3] , \dc32_fifo_data_out[2] , \dc32_fifo_data_out[1] , 
            DEBUG_5_c_0, DEBUG_2_c, sc32_fifo_read_enable, n5367, n5366, 
            n5365, n5364, n5363, n5362, n5361, n5360, n5359, n5358, 
            n5357, n5356, n5355, n5354, n5353, n5352, n5351, n5350, 
            n5349, n5348, n5347, n5346, n5345, n5344, n5343, n5342, 
            n5341, n5340, n5339, n5338, n5337) /* synthesis syn_module_defined=1 */ ;
    output DEBUG_9_c_0;
    input SLM_CLK_c;
    input \dc32_fifo_data_out[31] ;
    input \dc32_fifo_data_out[30] ;
    input \dc32_fifo_data_out[29] ;
    input \dc32_fifo_data_out[28] ;
    input \dc32_fifo_data_out[27] ;
    input \dc32_fifo_data_out[26] ;
    input \dc32_fifo_data_out[25] ;
    input \dc32_fifo_data_out[24] ;
    input \dc32_fifo_data_out[23] ;
    output sc32_fifo_almost_empty;
    input reset_all;
    input \dc32_fifo_data_out[22] ;
    input \dc32_fifo_data_out[21] ;
    input \dc32_fifo_data_out[20] ;
    input \dc32_fifo_data_out[19] ;
    input \dc32_fifo_data_out[18] ;
    input \dc32_fifo_data_out[17] ;
    input \dc32_fifo_data_out[16] ;
    input \dc32_fifo_data_out[15] ;
    input \dc32_fifo_data_out[14] ;
    input \dc32_fifo_data_out[13] ;
    input \dc32_fifo_data_out[12] ;
    input \dc32_fifo_data_out[11] ;
    input \dc32_fifo_data_out[10] ;
    input \dc32_fifo_data_out[9] ;
    input \dc32_fifo_data_out[8] ;
    input \dc32_fifo_data_out[7] ;
    input \dc32_fifo_data_out[6] ;
    input GND_net;
    input \dc32_fifo_data_out[5] ;
    input \dc32_fifo_data_out[4] ;
    input \dc32_fifo_data_out[3] ;
    input \dc32_fifo_data_out[2] ;
    input \dc32_fifo_data_out[1] ;
    input DEBUG_5_c_0;
    input DEBUG_2_c;
    input sc32_fifo_read_enable;
    output n5367;
    output n5366;
    output n5365;
    output n5364;
    output n5363;
    output n5362;
    output n5361;
    output n5360;
    output n5359;
    output n5358;
    output n5357;
    output n5356;
    output n5355;
    output n5354;
    output n5353;
    output n5352;
    output n5351;
    output n5350;
    output n5349;
    output n5348;
    output n5347;
    output n5346;
    output n5345;
    output n5344;
    output n5343;
    output n5342;
    output n5341;
    output n5340;
    output n5339;
    output n5338;
    output n5337;
>>>>>>> Stashed changes
>>>>>>> master
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
<<<<<<< HEAD
    fifo_sc_32_lut_gen_ipgen_lscc_fifo_renamed_due_excessive_length_2 lscc_fifo_inst (.SLM_CLK_c(SLM_CLK_c), 
            .sc32_fifo_almost_empty(sc32_fifo_almost_empty), .reset_all(reset_all), 
            .GND_net(GND_net), .dc32_fifo_read_enable(dc32_fifo_read_enable), 
            .sc32_fifo_read_enable(sc32_fifo_read_enable)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_sc_32_lut_gen.v(45[37] 59[45])
=======
<<<<<<< Updated upstream
    SB_PLL40_CORE pll_config (.REFERENCECLK(ICE_SYSCLK_c), .PLLOUTGLOBAL(pll_clk_unbuf), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=222, LSE_RLINE=228 */ ;   // src/top.v(222[7] 228[3])
    defparam pll_config.FEEDBACK_PATH = "SIMPLE";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll_config.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll_config.FDA_FEEDBACK = 0;
    defparam pll_config.FDA_RELATIVE = 0;
    defparam pll_config.PLLOUT_SELECT = "GENCLK";
    defparam pll_config.DIVR = 4'b0001;
    defparam pll_config.DIVF = 7'b1010010;
    defparam pll_config.DIVQ = 3'b100;
    defparam pll_config.FILTER_RANGE = 3'b001;
    defparam pll_config.ENABLE_ICEGATE = 1'b0;
    defparam pll_config.TEST_MODE = 1'b0;
    defparam pll_config.EXTERNAL_DIVIDE_FACTOR = 1;
=======
    fifo_sc_32_lut_gen_ipgen_lscc_fifo_renamed_due_excessive_length_2 lscc_fifo_inst (.DEBUG_9_c_0(DEBUG_9_c_0), 
            .SLM_CLK_c(SLM_CLK_c), .\dc32_fifo_data_out[31] (\dc32_fifo_data_out[31] ), 
            .\dc32_fifo_data_out[30] (\dc32_fifo_data_out[30] ), .\dc32_fifo_data_out[29] (\dc32_fifo_data_out[29] ), 
            .\dc32_fifo_data_out[28] (\dc32_fifo_data_out[28] ), .\dc32_fifo_data_out[27] (\dc32_fifo_data_out[27] ), 
            .\dc32_fifo_data_out[26] (\dc32_fifo_data_out[26] ), .\dc32_fifo_data_out[25] (\dc32_fifo_data_out[25] ), 
            .\dc32_fifo_data_out[24] (\dc32_fifo_data_out[24] ), .\dc32_fifo_data_out[23] (\dc32_fifo_data_out[23] ), 
            .sc32_fifo_almost_empty(sc32_fifo_almost_empty), .reset_all(reset_all), 
            .\dc32_fifo_data_out[22] (\dc32_fifo_data_out[22] ), .\dc32_fifo_data_out[21] (\dc32_fifo_data_out[21] ), 
            .\dc32_fifo_data_out[20] (\dc32_fifo_data_out[20] ), .\dc32_fifo_data_out[19] (\dc32_fifo_data_out[19] ), 
            .\dc32_fifo_data_out[18] (\dc32_fifo_data_out[18] ), .\dc32_fifo_data_out[17] (\dc32_fifo_data_out[17] ), 
            .\dc32_fifo_data_out[16] (\dc32_fifo_data_out[16] ), .\dc32_fifo_data_out[15] (\dc32_fifo_data_out[15] ), 
            .\dc32_fifo_data_out[14] (\dc32_fifo_data_out[14] ), .\dc32_fifo_data_out[13] (\dc32_fifo_data_out[13] ), 
            .\dc32_fifo_data_out[12] (\dc32_fifo_data_out[12] ), .\dc32_fifo_data_out[11] (\dc32_fifo_data_out[11] ), 
            .\dc32_fifo_data_out[10] (\dc32_fifo_data_out[10] ), .\dc32_fifo_data_out[9] (\dc32_fifo_data_out[9] ), 
            .\dc32_fifo_data_out[8] (\dc32_fifo_data_out[8] ), .\dc32_fifo_data_out[7] (\dc32_fifo_data_out[7] ), 
            .\dc32_fifo_data_out[6] (\dc32_fifo_data_out[6] ), .GND_net(GND_net), 
            .\dc32_fifo_data_out[5] (\dc32_fifo_data_out[5] ), .\dc32_fifo_data_out[4] (\dc32_fifo_data_out[4] ), 
            .\dc32_fifo_data_out[3] (\dc32_fifo_data_out[3] ), .\dc32_fifo_data_out[2] (\dc32_fifo_data_out[2] ), 
            .\dc32_fifo_data_out[1] (\dc32_fifo_data_out[1] ), .DEBUG_5_c_0(DEBUG_5_c_0), 
            .DEBUG_2_c(DEBUG_2_c), .sc32_fifo_read_enable(sc32_fifo_read_enable), 
            .n5367(n5367), .n5366(n5366), .n5365(n5365), .n5364(n5364), 
            .n5363(n5363), .n5362(n5362), .n5361(n5361), .n5360(n5360), 
            .n5359(n5359), .n5358(n5358), .n5357(n5357), .n5356(n5356), 
            .n5355(n5355), .n5354(n5354), .n5353(n5353), .n5352(n5352), 
            .n5351(n5351), .n5350(n5350), .n5349(n5349), .n5348(n5348), 
            .n5347(n5347), .n5346(n5346), .n5345(n5345), .n5344(n5344), 
            .n5343(n5343), .n5342(n5342), .n5341(n5341), .n5340(n5340), 
            .n5339(n5339), .n5338(n5338), .n5337(n5337)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_sc_32_lut_gen.v(45[37] 59[45])
>>>>>>> Stashed changes
>>>>>>> master
    
endmodule
//
// Verilog Description of module fifo_sc_32_lut_gen_ipgen_lscc_fifo_renamed_due_excessive_length_2
//

<<<<<<< HEAD
module fifo_sc_32_lut_gen_ipgen_lscc_fifo_renamed_due_excessive_length_2 (SLM_CLK_c, 
            sc32_fifo_almost_empty, reset_all, GND_net, dc32_fifo_read_enable, 
            sc32_fifo_read_enable) /* synthesis syn_module_defined=1 */ ;
=======
<<<<<<< Updated upstream
module \uart_rx(CLKS_PER_BIT=20)  (r_SM_Main, SLM_CLK_c, r_Rx_Data, GND_net, 
            n4, n4_adj_1, n6105, pc_data_rx, n10406, VCC_net, debug_led3, 
            n7473, n6082, n6081, n6079, n6078, n6077, n6075, n6074, 
            \r_SM_Main_2__N_765[2] , n4_adj_2, n10345, UART_RX_c, n4248, 
            n4253) /* synthesis syn_module_defined=1 */ ;
    output [2:0]r_SM_Main;
>>>>>>> master
    input SLM_CLK_c;
    output sc32_fifo_almost_empty;
    input reset_all;
    input GND_net;
    input dc32_fifo_read_enable;
    input sc32_fifo_read_enable;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire full_ext_r_N_793, full_r, empty_ext_r_N_795, empty_r;
    wire [3:0]wr_addr_r_3__N_689;
    wire [3:0]\MISC.wr_flag_addr_r ;   // src/fifo_sc_32_lut_gen.v(261[56:70])
    wire [3:0]wr_addr_p1_r_3__N_693;
    wire [3:0]\MISC.wr_flag_addr_p1_r ;   // src/fifo_sc_32_lut_gen.v(262[56:73])
    wire [3:0]rd_addr_r_3__N_707;
    wire [3:0]\MISC.rd_flag_addr_r ;   // src/fifo_sc_32_lut_gen.v(263[56:70])
    wire [3:0]rd_addr_p1_r_3__N_711;
    wire [3:0]\MISC.rd_flag_addr_p1_r ;   // src/fifo_sc_32_lut_gen.v(264[56:73])
    
    wire \MISC.AEmpty.almost_empty_nxt_w ;
    wire [3:0]n2649;
    
    wire n3293, n2, n4;
    wire [3:0]rd_addr_r;   // src/fifo_sc_32_lut_gen.v(123[48:57])
    wire [3:0]rd_addr_p1_r;   // src/fifo_sc_32_lut_gen.v(124[48:60])
    
    wire n3799, n3291, n3300, n2249, n10465, n4_adj_1366, n10466, 
        n6;
    wire [3:0]rd_addr_nxt_w;   // src/fifo_sc_32_lut_gen.v(133[28:41])
    wire [3:0]wr_addr_nxt_w;   // src/fifo_sc_32_lut_gen.v(130[28:41])
    wire [3:0]wr_addr_r;   // src/fifo_sc_32_lut_gen.v(117[48:57])
    
    wire n11149, n11223, wr_addr_nxt_w_3__N_728, n11269, full_nxt_w_N_811, 
        empty_nxt_w_N_822, rd_addr_nxt_w_3__N_732, n4_adj_1367;
    wire [3:0]wr_addr_p1_r;   // src/fifo_sc_32_lut_gen.v(118[48:60])
    
    wire n6_adj_1368, n11161, full_nxt_w_N_796, n11151;
    wire [2:0]rd_cmpaddr_p1_r_2__N_725;
    wire [2:0]rd_cmpaddr_r_2__N_719;
    wire [3:0]wr_addr_p1cmp_r_3__N_697;
    wire [2:0]wr_cmpaddr_p1_r_2__N_704;
    wire [2:0]wr_cmpaddr_r_2__N_698;
    
    wire n2965, n2994;
    
    SB_DFF full_r_122 (.Q(full_r), .C(SLM_CLK_c), .D(full_ext_r_N_793));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF empty_r_125 (.Q(empty_r), .C(SLM_CLK_c), .D(empty_ext_r_N_795));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF \MISC.wr_flag_addr_r_i0  (.Q(\MISC.wr_flag_addr_r [0]), .C(SLM_CLK_c), 
           .D(wr_addr_r_3__N_689[0]));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_DFF \MISC.wr_flag_addr_p1_r_i0  (.Q(\MISC.wr_flag_addr_p1_r [0]), .C(SLM_CLK_c), 
           .D(wr_addr_p1_r_3__N_693[0]));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_DFF \MISC.rd_flag_addr_r_i0  (.Q(\MISC.rd_flag_addr_r [0]), .C(SLM_CLK_c), 
           .D(rd_addr_r_3__N_707[0]));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_DFF \MISC.rd_flag_addr_p1_r_i0  (.Q(\MISC.rd_flag_addr_p1_r [0]), .C(SLM_CLK_c), 
           .D(rd_addr_p1_r_3__N_711[0]));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_DFFSS \MISC.AEmpty.almost_empty_ext_r_147  (.Q(sc32_fifo_almost_empty), 
            .C(SLM_CLK_c), .D(\MISC.AEmpty.almost_empty_nxt_w ), .S(reset_all));   // src/fifo_sc_32_lut_gen.v(403[33] 415[36])
    SB_LUT4 i1661_3_lut (.I0(n2649[1]), .I1(n3293), .I2(n2), .I3(GND_net), 
            .O(n4));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i1661_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i2353_3_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1_r[2]), .I2(n3799), 
            .I3(GND_net), .O(n3291));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i2353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2355_3_lut (.I0(rd_addr_r[1]), .I1(rd_addr_p1_r[1]), .I2(n3799), 
            .I3(GND_net), .O(n3293));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i2355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2037_3_lut (.I0(\MISC.rd_flag_addr_r [0]), .I1(\MISC.rd_flag_addr_p1_r [0]), 
            .I2(n3799), .I3(GND_net), .O(n3300));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i2037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1653_4_lut (.I0(\MISC.wr_flag_addr_r [0]), .I1(n3300), .I2(\MISC.wr_flag_addr_p1_r [0]), 
            .I3(n2249), .O(n2));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i1653_4_lut.LUT_INIT = 16'hf3bb;
    SB_LUT4 i2_3_lut (.I0(n2), .I1(n3293), .I2(n2649[1]), .I3(GND_net), 
            .O(n10465));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut (.I0(\MISC.rd_flag_addr_r [3]), .I1(n2649[3]), .I2(rd_addr_p1_r[3]), 
            .I3(n3799), .O(n4_adj_1366));
    defparam i1_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i2_3_lut_adj_42 (.I0(n4), .I1(n3291), .I2(n2649[2]), .I3(GND_net), 
            .O(n10466));
    defparam i2_3_lut_adj_42.LUT_INIT = 16'h9696;
    SB_LUT4 i1668_3_lut (.I0(n2649[2]), .I1(n3291), .I2(n4), .I3(GND_net), 
            .O(n6));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i1668_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i2_4_lut (.I0(n6), .I1(n10466), .I2(n4_adj_1366), .I3(n10465), 
            .O(\MISC.AEmpty.almost_empty_nxt_w ));
    defparam i2_4_lut.LUT_INIT = 16'h4800;
    SB_LUT4 i6375_2_lut (.I0(rd_addr_nxt_w[0]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(rd_addr_p1_r_3__N_711[0]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6375_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i6374_2_lut (.I0(rd_addr_nxt_w[0]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(rd_addr_r_3__N_707[0]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6374_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6372_2_lut (.I0(wr_addr_nxt_w[0]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(wr_addr_p1_r_3__N_693[0]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6372_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i6365_2_lut (.I0(wr_addr_nxt_w[0]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(wr_addr_r_3__N_689[0]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6365_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i9573_4_lut (.I0(rd_addr_p1_r[2]), .I1(rd_addr_p1_r[3]), .I2(wr_addr_r[2]), 
            .I3(\MISC.wr_flag_addr_r [3]), .O(n11149));
    defparam i9573_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i9646_3_lut (.I0(\MISC.rd_flag_addr_p1_r [0]), .I1(n11149), 
            .I2(\MISC.wr_flag_addr_r [0]), .I3(GND_net), .O(n11223));
    defparam i9646_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 i9691_4_lut (.I0(rd_addr_p1_r[1]), .I1(n11223), .I2(wr_addr_nxt_w_3__N_728), 
            .I3(wr_addr_r[1]), .O(n11269));
    defparam i9691_4_lut.LUT_INIT = 16'hfdfe;
    SB_LUT4 i2_3_lut_adj_43 (.I0(empty_r), .I1(dc32_fifo_read_enable), .I2(full_nxt_w_N_811), 
            .I3(GND_net), .O(empty_nxt_w_N_822));
    defparam i2_3_lut_adj_43.LUT_INIT = 16'h0202;
    SB_LUT4 i1_4_lut_adj_44 (.I0(reset_all), .I1(rd_addr_nxt_w_3__N_732), 
            .I2(empty_nxt_w_N_822), .I3(n11269), .O(empty_ext_r_N_795));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i1_4_lut_adj_44.LUT_INIT = 16'hfafe;
    SB_LUT4 i1_4_lut_adj_45 (.I0(wr_addr_r[2]), .I1(\MISC.wr_flag_addr_r [0]), 
            .I2(rd_addr_r[2]), .I3(\MISC.rd_flag_addr_r [0]), .O(n4_adj_1367));   // src/fifo_sc_32_lut_gen.v(136[186:216])
    defparam i1_4_lut_adj_45.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_3_lut_adj_46 (.I0(wr_addr_r[1]), .I1(n4_adj_1367), .I2(rd_addr_r[1]), 
            .I3(GND_net), .O(full_nxt_w_N_811));   // src/fifo_sc_32_lut_gen.v(136[186:216])
    defparam i2_3_lut_adj_46.LUT_INIT = 16'hdede;
    SB_LUT4 wr_en_i_I_0_167_2_lut (.I0(dc32_fifo_read_enable), .I1(full_r), 
            .I2(GND_net), .I3(GND_net), .O(wr_addr_nxt_w_3__N_728));   // src/fifo_sc_32_lut_gen.v(130[45:66])
    defparam wr_en_i_I_0_167_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 rd_en_i_I_0_165_2_lut (.I0(sc32_fifo_read_enable), .I1(empty_r), 
            .I2(GND_net), .I3(GND_net), .O(rd_addr_nxt_w_3__N_732));   // src/fifo_sc_32_lut_gen.v(133[45:67])
    defparam rd_en_i_I_0_165_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_4_lut_adj_47 (.I0(wr_addr_p1_r[3]), .I1(wr_addr_p1_r[1]), 
            .I2(\MISC.rd_flag_addr_r [3]), .I3(rd_addr_r[1]), .O(n6_adj_1368));
    defparam i2_4_lut_adj_47.LUT_INIT = 16'h4812;
    SB_LUT4 i9585_4_lut (.I0(\MISC.wr_flag_addr_p1_r [0]), .I1(wr_addr_p1_r[2]), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(rd_addr_r[2]), .O(n11161));
    defparam i9585_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_3_lut_adj_48 (.I0(n11161), .I1(n2249), .I2(n6_adj_1368), 
            .I3(GND_net), .O(full_nxt_w_N_796));
    defparam i2_3_lut_adj_48.LUT_INIT = 16'h4040;
    SB_LUT4 i6370_4_lut (.I0(full_nxt_w_N_796), .I1(reset_all), .I2(full_r), 
            .I3(n11151), .O(full_ext_r_N_793));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6370_4_lut.LUT_INIT = 16'h2232;
    SB_DFF \MISC.rd_flag_addr_r_i3  (.Q(\MISC.rd_flag_addr_r [3]), .C(SLM_CLK_c), 
           .D(rd_addr_r_3__N_707[3]));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_DFF \MISC.wr_flag_addr_r_i3  (.Q(\MISC.wr_flag_addr_r [3]), .C(SLM_CLK_c), 
           .D(wr_addr_r_3__N_689[3]));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_DFF rd_addr_p1_r_i3 (.Q(rd_addr_p1_r[3]), .C(SLM_CLK_c), .D(rd_addr_p1_r_3__N_711[3]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF rd_addr_p1_r_i2 (.Q(rd_addr_p1_r[2]), .C(SLM_CLK_c), .D(rd_cmpaddr_p1_r_2__N_725[2]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF rd_addr_p1_r_i1 (.Q(rd_addr_p1_r[1]), .C(SLM_CLK_c), .D(rd_cmpaddr_p1_r_2__N_725[1]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF rd_addr_r_i2 (.Q(rd_addr_r[2]), .C(SLM_CLK_c), .D(rd_cmpaddr_r_2__N_719[2]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF rd_addr_r_i1 (.Q(rd_addr_r[1]), .C(SLM_CLK_c), .D(rd_cmpaddr_r_2__N_719[1]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF wr_addr_p1_r_i3 (.Q(wr_addr_p1_r[3]), .C(SLM_CLK_c), .D(wr_addr_p1cmp_r_3__N_697[3]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF wr_addr_p1_r_i2 (.Q(wr_addr_p1_r[2]), .C(SLM_CLK_c), .D(wr_cmpaddr_p1_r_2__N_704[2]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF wr_addr_p1_r_i1 (.Q(wr_addr_p1_r[1]), .C(SLM_CLK_c), .D(wr_cmpaddr_p1_r_2__N_704[1]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF wr_addr_r_i2 (.Q(wr_addr_r[2]), .C(SLM_CLK_c), .D(wr_cmpaddr_r_2__N_698[2]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF wr_addr_r_i1 (.Q(wr_addr_r[1]), .C(SLM_CLK_c), .D(wr_cmpaddr_r_2__N_698[1]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_LUT4 i6437_2_lut (.I0(wr_addr_nxt_w[1]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(wr_cmpaddr_r_2__N_698[1]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6437_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6436_2_lut (.I0(wr_addr_nxt_w[2]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(wr_cmpaddr_r_2__N_698[2]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6436_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6435_3_lut (.I0(wr_addr_nxt_w[1]), .I1(reset_all), .I2(wr_addr_nxt_w[0]), 
            .I3(GND_net), .O(wr_cmpaddr_p1_r_2__N_704[1]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6435_3_lut.LUT_INIT = 16'h1212;
    SB_LUT4 i1556_2_lut (.I0(wr_addr_nxt_w[1]), .I1(wr_addr_nxt_w[0]), .I2(GND_net), 
            .I3(GND_net), .O(n2965));   // src/fifo_sc_32_lut_gen.v(131[47:69])
    defparam i1556_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6373_4_lut (.I0(wr_addr_nxt_w[3]), .I1(reset_all), .I2(wr_addr_nxt_w[2]), 
            .I3(n2965), .O(wr_addr_p1cmp_r_3__N_697[3]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6373_4_lut.LUT_INIT = 16'h1222;
    SB_LUT4 i6431_2_lut (.I0(rd_addr_nxt_w[1]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(rd_cmpaddr_r_2__N_719[1]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6431_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6430_2_lut (.I0(rd_addr_nxt_w[2]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(rd_cmpaddr_r_2__N_719[2]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6430_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6429_3_lut (.I0(rd_addr_nxt_w[1]), .I1(reset_all), .I2(rd_addr_nxt_w[0]), 
            .I3(GND_net), .O(rd_cmpaddr_p1_r_2__N_725[1]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6429_3_lut.LUT_INIT = 16'h1212;
    SB_LUT4 i2350_3_lut_4_lut_4_lut (.I0(dc32_fifo_read_enable), .I1(full_r), 
            .I2(sc32_fifo_read_enable), .I3(empty_r), .O(n3799));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i2350_3_lut_4_lut_4_lut.LUT_INIT = 16'h00d0;
    SB_LUT4 i1585_2_lut (.I0(rd_addr_nxt_w[1]), .I1(rd_addr_nxt_w[0]), .I2(GND_net), 
            .I3(GND_net), .O(n2994));   // src/fifo_sc_32_lut_gen.v(134[47:69])
    defparam i1585_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6432_4_lut (.I0(rd_addr_nxt_w[3]), .I1(reset_all), .I2(rd_addr_nxt_w[2]), 
            .I3(n2994), .O(rd_addr_p1_r_3__N_711[3]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6432_4_lut.LUT_INIT = 16'h1222;
    SB_LUT4 i6438_2_lut (.I0(wr_addr_nxt_w[3]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(wr_addr_r_3__N_689[3]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6438_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6433_2_lut (.I0(rd_addr_nxt_w[3]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(rd_addr_r_3__N_707[3]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6433_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 rd_addr_r_3__I_0_i4_3_lut_4_lut (.I0(\MISC.rd_flag_addr_r [3]), 
            .I1(rd_addr_p1_r[3]), .I2(sc32_fifo_read_enable), .I3(empty_r), 
            .O(rd_addr_nxt_w[3]));   // src/fifo_sc_32_lut_gen.v(133[44:95])
    defparam rd_addr_r_3__I_0_i4_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 wr_addr_r_3__I_0_i4_3_lut_4_lut (.I0(\MISC.wr_flag_addr_r [3]), 
            .I1(wr_addr_p1_r[3]), .I2(dc32_fifo_read_enable), .I3(full_r), 
            .O(wr_addr_nxt_w[3]));   // src/fifo_sc_32_lut_gen.v(130[44:94])
    defparam wr_addr_r_3__I_0_i4_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 rd_addr_r_3__I_0_i3_3_lut_4_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1_r[2]), 
            .I2(sc32_fifo_read_enable), .I3(empty_r), .O(rd_addr_nxt_w[2]));   // src/fifo_sc_32_lut_gen.v(133[44:95])
    defparam rd_addr_r_3__I_0_i3_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 rd_addr_r_3__I_0_i2_3_lut_4_lut (.I0(rd_addr_r[1]), .I1(rd_addr_p1_r[1]), 
            .I2(sc32_fifo_read_enable), .I3(empty_r), .O(rd_addr_nxt_w[1]));   // src/fifo_sc_32_lut_gen.v(133[44:95])
    defparam rd_addr_r_3__I_0_i2_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i6428_3_lut_4_lut (.I0(rd_addr_nxt_w[2]), .I1(reset_all), .I2(rd_addr_nxt_w[1]), 
            .I3(rd_addr_nxt_w[0]), .O(rd_cmpaddr_p1_r_2__N_725[2]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6428_3_lut_4_lut.LUT_INIT = 16'h1222;
    SB_LUT4 wr_addr_r_3__I_0_i3_3_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_r[2]), 
            .I2(dc32_fifo_read_enable), .I3(full_r), .O(wr_addr_nxt_w[2]));   // src/fifo_sc_32_lut_gen.v(130[44:94])
    defparam wr_addr_r_3__I_0_i3_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 wr_addr_r_3__I_0_i2_3_lut_4_lut (.I0(wr_addr_r[1]), .I1(wr_addr_p1_r[1]), 
            .I2(dc32_fifo_read_enable), .I3(full_r), .O(wr_addr_nxt_w[1]));   // src/fifo_sc_32_lut_gen.v(130[44:94])
    defparam wr_addr_r_3__I_0_i2_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i6434_3_lut_4_lut (.I0(wr_addr_nxt_w[2]), .I1(reset_all), .I2(wr_addr_nxt_w[1]), 
            .I3(wr_addr_nxt_w[0]), .O(wr_cmpaddr_p1_r_2__N_704[2]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i6434_3_lut_4_lut.LUT_INIT = 16'h1222;
    SB_LUT4 i9575_2_lut_4_lut (.I0(sc32_fifo_read_enable), .I1(wr_addr_r[1]), 
            .I2(n4_adj_1367), .I3(rd_addr_r[1]), .O(n11151));
    defparam i9575_2_lut_4_lut.LUT_INIT = 16'hfbfe;
    SB_LUT4 i1077_2_lut_4_lut (.I0(sc32_fifo_read_enable), .I1(empty_r), 
            .I2(dc32_fifo_read_enable), .I3(full_r), .O(n2249));   // src/fifo_sc_32_lut_gen.v(270[46:60])
    defparam i1077_2_lut_4_lut.LUT_INIT = 16'h00d0;
    SB_LUT4 wr_addr_r_3__I_0_i1_3_lut_4_lut (.I0(\MISC.wr_flag_addr_r [0]), 
            .I1(\MISC.wr_flag_addr_p1_r [0]), .I2(dc32_fifo_read_enable), 
            .I3(full_r), .O(wr_addr_nxt_w[0]));   // src/fifo_sc_32_lut_gen.v(130[44:94])
    defparam wr_addr_r_3__I_0_i1_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 rd_addr_r_3__I_0_i1_3_lut_4_lut (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\MISC.rd_flag_addr_p1_r [0]), .I2(sc32_fifo_read_enable), 
            .I3(empty_r), .O(rd_addr_nxt_w[0]));   // src/fifo_sc_32_lut_gen.v(133[44:95])
    defparam rd_addr_r_3__I_0_i1_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 mux_1336_i4_3_lut_4_lut (.I0(\MISC.wr_flag_addr_r [3]), .I1(wr_addr_p1_r[3]), 
            .I2(rd_addr_nxt_w_3__N_732), .I3(wr_addr_nxt_w_3__N_728), .O(n2649[3]));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam mux_1336_i4_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_1336_i2_3_lut_4_lut (.I0(wr_addr_r[1]), .I1(wr_addr_p1_r[1]), 
            .I2(rd_addr_nxt_w_3__N_732), .I3(wr_addr_nxt_w_3__N_728), .O(n2649[1]));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam mux_1336_i2_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_1336_i3_3_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_r[2]), 
            .I2(rd_addr_nxt_w_3__N_732), .I3(wr_addr_nxt_w_3__N_728), .O(n2649[2]));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam mux_1336_i3_3_lut_4_lut.LUT_INIT = 16'hacaa;
    
endmodule
//
// Verilog Description of module FIFO_Quad_Word
//

module FIFO_Quad_Word (rd_addr_r, SLM_CLK_c, reset_all_w, \mem_LUT.data_raw_r[0] , 
            wr_addr_r, fifo_write_cmd, is_tx_fifo_full_flag, wr_fifo_en_w, 
            GND_net, n2704, \wr_addr_p1_w[2] , n1, n10381, \mem_LUT.data_raw_r[7] , 
            \mem_LUT.data_raw_r[6] , \mem_LUT.data_raw_r[5] , \mem_LUT.data_raw_r[4] , 
            \mem_LUT.data_raw_r[3] , \mem_LUT.data_raw_r[2] , \mem_LUT.data_raw_r[1] , 
            rx_buf_byte, n5734, \fifo_temp_output[1] , n10640, VCC_net, 
            n5738, \fifo_temp_output[2] , n5633, rd_fifo_en_prev_r, 
            fifo_read_cmd, is_fifo_empty_flag, empty_o_N_1333, n11046, 
            n5741, \fifo_temp_output[3] , n5745, \fifo_temp_output[4] , 
            n5748, \fifo_temp_output[5] , n5812, \fifo_temp_output[0] , 
            n5755, \fifo_temp_output[6] , n5761, \fifo_temp_output[7] , 
            n5769, n5610, n5614, \rd_addr_p1_w[2] , n11863) /* synthesis syn_module_defined=1 */ ;
    output [2:0]rd_addr_r;
    input SLM_CLK_c;
    input reset_all_w;
    output \mem_LUT.data_raw_r[0] ;
    output [2:0]wr_addr_r;
    input fifo_write_cmd;
    output is_tx_fifo_full_flag;
    output wr_fifo_en_w;
    input GND_net;
    input n2704;
    output \wr_addr_p1_w[2] ;
    output n1;
    output n10381;
    output \mem_LUT.data_raw_r[7] ;
    output \mem_LUT.data_raw_r[6] ;
    output \mem_LUT.data_raw_r[5] ;
    output \mem_LUT.data_raw_r[4] ;
    output \mem_LUT.data_raw_r[3] ;
    output \mem_LUT.data_raw_r[2] ;
    output \mem_LUT.data_raw_r[1] ;
    input [7:0]rx_buf_byte;
    input n5734;
    output \fifo_temp_output[1] ;
    input n10640;
    input VCC_net;
    input n5738;
    output \fifo_temp_output[2] ;
    input n5633;
    output rd_fifo_en_prev_r;
    input fifo_read_cmd;
    output is_fifo_empty_flag;
    input empty_o_N_1333;
    input n11046;
    input n5741;
    output \fifo_temp_output[3] ;
    input n5745;
    output \fifo_temp_output[4] ;
    input n5748;
    output \fifo_temp_output[5] ;
    input n5812;
    output \fifo_temp_output[0] ;
    input n5755;
    output \fifo_temp_output[6] ;
    input n5761;
    output \fifo_temp_output[7] ;
<<<<<<< HEAD
    input n5769;
    input n5610;
    input n5614;
    output \rd_addr_p1_w[2] ;
    output n11863;
=======
    input n10786;
    output is_fifo_empty_flag;
    input n4919;
    input n4922;
    input fifo_write_cmd;
    output wr_fifo_en_w;
    input n4878;
    output rd_fifo_en_prev_r;
    input fifo_read_cmd;
=======
module fifo_sc_32_lut_gen_ipgen_lscc_fifo_renamed_due_excessive_length_2 (DEBUG_9_c_0, 
            SLM_CLK_c, \dc32_fifo_data_out[31] , \dc32_fifo_data_out[30] , 
            \dc32_fifo_data_out[29] , \dc32_fifo_data_out[28] , \dc32_fifo_data_out[27] , 
            \dc32_fifo_data_out[26] , \dc32_fifo_data_out[25] , \dc32_fifo_data_out[24] , 
            \dc32_fifo_data_out[23] , sc32_fifo_almost_empty, reset_all, 
            \dc32_fifo_data_out[22] , \dc32_fifo_data_out[21] , \dc32_fifo_data_out[20] , 
            \dc32_fifo_data_out[19] , \dc32_fifo_data_out[18] , \dc32_fifo_data_out[17] , 
            \dc32_fifo_data_out[16] , \dc32_fifo_data_out[15] , \dc32_fifo_data_out[14] , 
            \dc32_fifo_data_out[13] , \dc32_fifo_data_out[12] , \dc32_fifo_data_out[11] , 
            \dc32_fifo_data_out[10] , \dc32_fifo_data_out[9] , \dc32_fifo_data_out[8] , 
            \dc32_fifo_data_out[7] , \dc32_fifo_data_out[6] , GND_net, 
            \dc32_fifo_data_out[5] , \dc32_fifo_data_out[4] , \dc32_fifo_data_out[3] , 
            \dc32_fifo_data_out[2] , \dc32_fifo_data_out[1] , DEBUG_5_c_0, 
            DEBUG_2_c, sc32_fifo_read_enable, n5367, n5366, n5365, 
            n5364, n5363, n5362, n5361, n5360, n5359, n5358, n5357, 
            n5356, n5355, n5354, n5353, n5352, n5351, n5350, n5349, 
            n5348, n5347, n5346, n5345, n5344, n5343, n5342, n5341, 
            n5340, n5339, n5338, n5337) /* synthesis syn_module_defined=1 */ ;
    output DEBUG_9_c_0;
    input SLM_CLK_c;
    input \dc32_fifo_data_out[31] ;
    input \dc32_fifo_data_out[30] ;
    input \dc32_fifo_data_out[29] ;
    input \dc32_fifo_data_out[28] ;
    input \dc32_fifo_data_out[27] ;
    input \dc32_fifo_data_out[26] ;
    input \dc32_fifo_data_out[25] ;
    input \dc32_fifo_data_out[24] ;
    input \dc32_fifo_data_out[23] ;
    output sc32_fifo_almost_empty;
    input reset_all;
    input \dc32_fifo_data_out[22] ;
    input \dc32_fifo_data_out[21] ;
    input \dc32_fifo_data_out[20] ;
    input \dc32_fifo_data_out[19] ;
    input \dc32_fifo_data_out[18] ;
    input \dc32_fifo_data_out[17] ;
    input \dc32_fifo_data_out[16] ;
    input \dc32_fifo_data_out[15] ;
    input \dc32_fifo_data_out[14] ;
    input \dc32_fifo_data_out[13] ;
    input \dc32_fifo_data_out[12] ;
    input \dc32_fifo_data_out[11] ;
    input \dc32_fifo_data_out[10] ;
    input \dc32_fifo_data_out[9] ;
    input \dc32_fifo_data_out[8] ;
    input \dc32_fifo_data_out[7] ;
    input \dc32_fifo_data_out[6] ;
    input GND_net;
    input \dc32_fifo_data_out[5] ;
    input \dc32_fifo_data_out[4] ;
    input \dc32_fifo_data_out[3] ;
    input \dc32_fifo_data_out[2] ;
    input \dc32_fifo_data_out[1] ;
    input DEBUG_5_c_0;
    input DEBUG_2_c;
    input sc32_fifo_read_enable;
    output n5367;
    output n5366;
    output n5365;
    output n5364;
    output n5363;
    output n5362;
    output n5361;
    output n5360;
    output n5359;
    output n5358;
    output n5357;
    output n5356;
    output n5355;
    output n5354;
    output n5353;
    output n5352;
    output n5351;
    output n5350;
    output n5349;
    output n5348;
    output n5347;
    output n5346;
    output n5345;
    output n5344;
    output n5343;
    output n5342;
    output n5341;
    output n5340;
    output n5339;
    output n5338;
    output n5337;
>>>>>>> master
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [3:0]\MISC.rd_flag_addr_r ;   // src/fifo_sc_32_lut_gen.v(263[56:70])
    
    wire \mem_REG.mem_2_28 , \mem_REG.mem_3_28 ;
    wire [3:0]rd_addr_r;   // src/fifo_sc_32_lut_gen.v(123[48:57])
    
    wire n15781, \mem_REG.mem_1_28 , \mem_REG.mem_0_28 , n15784, \mem_REG.mem_2_13 , 
        \mem_REG.mem_3_13 , n14635;
    wire [31:0]rd_data_o_31__N_759;
    
<<<<<<< HEAD
    FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_3 lscc_fifo_inst (.rd_addr_r({rd_addr_r}), 
            .SLM_CLK_c(SLM_CLK_c), .reset_all_w(reset_all_w), .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r[0] ), 
            .wr_addr_r({wr_addr_r}), .fifo_write_cmd(fifo_write_cmd), .is_tx_fifo_full_flag(is_tx_fifo_full_flag), 
            .wr_fifo_en_w(wr_fifo_en_w), .GND_net(GND_net), .n2704(n2704), 
            .\wr_addr_p1_w[2] (\wr_addr_p1_w[2] ), .n1(n1), .n10381(n10381), 
            .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r[7] ), .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r[6] ), 
            .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r[5] ), .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r[4] ), 
            .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r[3] ), .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r[2] ), 
            .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r[1] ), .rx_buf_byte({rx_buf_byte}), 
            .n5734(n5734), .\fifo_temp_output[1] (\fifo_temp_output[1] ), 
            .n10640(n10640), .VCC_net(VCC_net), .n5738(n5738), .\fifo_temp_output[2] (\fifo_temp_output[2] ), 
            .n5633(n5633), .rd_fifo_en_prev_r(rd_fifo_en_prev_r), .fifo_read_cmd(fifo_read_cmd), 
            .is_fifo_empty_flag(is_fifo_empty_flag), .empty_o_N_1333(empty_o_N_1333), 
            .n11046(n11046), .n5741(n5741), .\fifo_temp_output[3] (\fifo_temp_output[3] ), 
            .n5745(n5745), .\fifo_temp_output[4] (\fifo_temp_output[4] ), 
            .n5748(n5748), .\fifo_temp_output[5] (\fifo_temp_output[5] ), 
            .n5812(n5812), .\fifo_temp_output[0] (\fifo_temp_output[0] ), 
            .n5755(n5755), .\fifo_temp_output[6] (\fifo_temp_output[6] ), 
            .n5761(n5761), .\fifo_temp_output[7] (\fifo_temp_output[7] ), 
            .n5769(n5769), .n5610(n5610), .n5614(n5614), .\rd_addr_p1_w[2] (\rd_addr_p1_w[2] ), 
            .n11863(n11863)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_quad_word_mod.v(20[37:380])
=======
    wire \MISC.rd_w , \mem_REG.mem_1_13 , \mem_REG.mem_0_13 , n14638, 
        \mem_REG.mem_6_28 , \mem_REG.mem_7_28 , n15739, \mem_REG.mem_5_28 , 
        \mem_REG.mem_4_28 , n15742, n13801, n13802, n15733, n13781, 
        n13780, n13807, n13808, n15727, n13784, n13783, n8;
    wire [3:0]wr_addr_r;   // src/fifo_sc_32_lut_gen.v(117[48:57])
    
    wire \mem_REG.mem_7_31 , n6877, \mem_REG.mem_7_30 , n6876, \mem_REG.mem_7_29 , 
        n6875;
    wire [3:0]wr_addr_r_3__N_690;
    wire [3:0]\MISC.wr_flag_addr_r ;   // src/fifo_sc_32_lut_gen.v(261[56:70])
    wire [3:0]wr_addr_p1_r_3__N_694;
    wire [3:0]\MISC.wr_flag_addr_p1_r ;   // src/fifo_sc_32_lut_gen.v(262[56:73])
    
    wire n6874;
    wire [3:0]rd_addr_r_3__N_708;
    
    wire \mem_REG.mem_7_27 , n6873, \mem_REG.mem_7_26 , n6872, \mem_REG.mem_7_25 , 
        n6871;
    wire [3:0]rd_addr_p1_r_3__N_712;
    wire [3:0]\MISC.rd_flag_addr_p1_r ;   // src/fifo_sc_32_lut_gen.v(264[56:73])
>>>>>>> Stashed changes
    
    wire \mem_REG.mem_7_24 , n6870, full_ext_r_N_794, \MISC.full_flag_r , 
        empty_ext_r_N_796, \MISC.empty_flag_r , \mem_REG.mem_7_23 , n6869, 
        \MISC.AEmpty.almost_empty_nxt_w , \mem_REG.mem_7_22 , n6868, \mem_REG.mem_7_21 , 
        n6867, \mem_REG.mem_7_20 , n6866, \mem_REG.mem_7_19 , n6865, 
        \mem_REG.mem_7_18 , n6864, \mem_REG.mem_7_17 , n6863, \mem_REG.mem_7_16 , 
        n6862, n13723, n13724, n15001, \mem_REG.mem_7_15 , n6861, 
        \mem_REG.mem_7_14 , n6860, \mem_REG.mem_7_13 , n6859, \mem_REG.mem_7_12 , 
        n6858, n13430, n13429, \mem_REG.mem_7_11 , n6857, \mem_REG.mem_7_10 , 
        n6856, \mem_REG.mem_7_9 , n6855, \mem_REG.mem_7_8 , n6854, 
        \mem_REG.mem_2_11 , \mem_REG.mem_3_11 , n15703, \mem_REG.mem_7_7 , 
        n6853, \mem_REG.mem_1_11 , \mem_REG.mem_0_11 , n15706, \mem_REG.mem_6_1 , 
        \mem_REG.mem_7_1 , n15697, \mem_REG.mem_5_1 , \mem_REG.mem_4_1 , 
        n15700, \mem_REG.mem_7_6 , n6852, \mem_REG.mem_0_8 , \mem_REG.mem_1_8 , 
        n13678, \mem_REG.mem_2_8 , \mem_REG.mem_3_8 , n13679, \mem_REG.mem_7_5 , 
        n6851, \mem_REG.mem_6_8 , n13709, \mem_REG.mem_4_8 , \mem_REG.mem_5_8 , 
        n13708, \mem_REG.mem_7_4 , n6850, \mem_REG.mem_7_3 , n6849, 
        n13732, n13733, n14983, \mem_REG.mem_7_2 , n6848, n6847, 
        n13151, n13150, \mem_REG.mem_7_0 , n6846, \mem_REG.mem_0_24 , 
        \mem_REG.mem_1_24 , n13720, \mem_REG.mem_2_24 , \mem_REG.mem_3_24 , 
        n13721, \mem_REG.mem_6_24 , n13727, \mem_REG.mem_4_24 , \mem_REG.mem_5_24 , 
        n13726, \mem_REG.mem_0_9 , \mem_REG.mem_1_9 , n13744, \mem_REG.mem_2_9 , 
        \mem_REG.mem_3_9 , n13745, \mem_REG.mem_6_9 , n13805, \mem_REG.mem_4_9 , 
        \mem_REG.mem_5_9 , n13804, \mem_REG.mem_0_2 , \mem_REG.mem_1_2 , 
        n13327, \mem_REG.mem_2_2 , \mem_REG.mem_3_2 , n13328, \mem_REG.mem_6_2 , 
        n13331, \mem_REG.mem_4_2 , \mem_REG.mem_5_2 , n13330, \mem_REG.mem_2_29 , 
        \mem_REG.mem_3_29 , n15679, \mem_REG.mem_1_29 , \mem_REG.mem_0_29 , 
        n15682, n13777, n13778, n15661, n13670, n13669, \mem_REG.mem_0_25 , 
        \mem_REG.mem_1_25 , n13753, \mem_REG.mem_2_25 , \mem_REG.mem_3_25 , 
        n13754, \mem_REG.mem_6_25 , n13673, \mem_REG.mem_4_25 , \mem_REG.mem_5_25 , 
        n13672, n6, \mem_REG.mem_6_31 , n6845, \mem_REG.mem_6_30 , 
        n6844, \mem_REG.mem_6_29 , n6843, n6842, \mem_REG.mem_6_27 , 
        n6841, \mem_REG.mem_6_26 , n6840, n6839, n6838, \mem_REG.mem_6_23 , 
        n6837, \mem_REG.mem_6_22 , n6836, \mem_REG.mem_6_21 , n6835, 
        \mem_REG.mem_6_20 , n6834, \mem_REG.mem_6_19 , n6833, \mem_REG.mem_6_18 , 
        n6832, \mem_REG.mem_6_17 , n6831, \mem_REG.mem_6_16 , n6830, 
        \mem_REG.mem_6_15 , n6829, \mem_REG.mem_6_14 , n6828, \mem_REG.mem_6_13 , 
        n6827, \mem_REG.mem_6_12 , n6826, \mem_REG.mem_6_11 , n6825, 
        \mem_REG.mem_6_10 , n6824, n6823, n6822, \mem_REG.mem_6_7 , 
        n6821, \mem_REG.mem_6_6 , n6820, \mem_REG.mem_6_5 , n6819, 
        \mem_REG.mem_6_4 , n6818, \mem_REG.mem_6_3 , n6817, n6816, 
        n6815, \mem_REG.mem_6_0 , n6814, n6813, \mem_REG.mem_5_31 , 
        n6812, \mem_REG.mem_5_30 , n6811, \mem_REG.mem_5_29 , n6810, 
        n6809, \mem_REG.mem_5_27 , n6808, \mem_REG.mem_5_26 , n6807, 
        n6806, n6805, \mem_REG.mem_5_23 , n6804, \mem_REG.mem_5_22 , 
        n6803, \mem_REG.mem_5_21 , n6802, \mem_REG.mem_5_20 , n6801, 
        \mem_REG.mem_5_19 , n6800, \mem_REG.mem_5_18 , n6799, \mem_REG.mem_5_17 , 
        n6798, \mem_REG.mem_5_16 , n6797, \mem_REG.mem_5_15 , n6796, 
        \mem_REG.mem_5_14 , n6795, \mem_REG.mem_5_13 , n6794, \mem_REG.mem_5_12 , 
        n6793, \mem_REG.mem_5_11 , n6792, \mem_REG.mem_5_10 , n6791, 
        n6790, n6789, \mem_REG.mem_5_7 , n6788, \mem_REG.mem_5_6 , 
        n6787, \mem_REG.mem_5_5 , n6786, \mem_REG.mem_5_4 , n6785, 
        \mem_REG.mem_5_3 , n6784, n6783, n6782, \mem_REG.mem_5_0 , 
        n6781, \mem_REG.mem_4_31 , n6780, \mem_REG.mem_4_30 , n6779, 
        \mem_REG.mem_4_29 , n6778, n6777, \mem_REG.mem_4_27 , n6776, 
        \mem_REG.mem_4_26 , n6775, n6774, n6773, \mem_REG.mem_4_23 , 
        n6772, \mem_REG.mem_4_22 , n6771, \mem_REG.mem_4_21 , n6770, 
        \mem_REG.mem_4_20 , n6769, \mem_REG.mem_4_19 , n6768, \mem_REG.mem_4_18 , 
        n6767, \mem_REG.mem_4_17 , n6766, \mem_REG.mem_4_16 , n6765, 
        \mem_REG.mem_4_15 , n6764, \mem_REG.mem_4_14 , n6763, \mem_REG.mem_4_13 , 
        n6762, \mem_REG.mem_4_12 , n6761, \mem_REG.mem_4_11 , n6760, 
        \mem_REG.mem_4_10 , n6759, n6758, n6757, \mem_REG.mem_4_7 , 
        n6756, \mem_REG.mem_4_6 , n6755, \mem_REG.mem_4_5 , n6754, 
        \mem_REG.mem_4_4 , n6753, \mem_REG.mem_4_3 , n6752, n6751, 
        n6750, \mem_REG.mem_4_0 , n6749, \mem_REG.mem_3_31 , n6748, 
        \mem_REG.mem_3_30 , n6747, n6746, n6745, \mem_REG.mem_3_27 , 
        n6744, \mem_REG.mem_3_26 , n6743, n6742, n6741, \mem_REG.mem_3_23 , 
        n6740, \mem_REG.mem_3_22 , n6739, \mem_REG.mem_3_21 , n6738, 
        \mem_REG.mem_3_20 , n6737, \mem_REG.mem_3_19 , n6736, \mem_REG.mem_3_18 , 
        n6735, \mem_REG.mem_3_17 , n6734, \mem_REG.mem_3_16 , n6733, 
        \mem_REG.mem_3_15 , n6732, \mem_REG.mem_3_14 , n6731, n6730, 
        \mem_REG.mem_3_12 , n6729, n6728, \mem_REG.mem_3_10 , n6727, 
        n6726, n6725, \mem_REG.mem_3_7 , n6724, \mem_REG.mem_3_6 , 
        n6723, \mem_REG.mem_3_5 , n6722, \mem_REG.mem_3_4 , n6721, 
        \mem_REG.mem_3_3 , n6720, n6719, \mem_REG.mem_3_1 , n6718, 
        \mem_REG.mem_3_0 , n6717, \mem_REG.mem_2_31 , n6716, \mem_REG.mem_2_30 , 
        n6715, n6714, n6713, \mem_REG.mem_2_27 , n6712, \mem_REG.mem_2_26 , 
        n6711, n6710, n6709, \mem_REG.mem_2_23 , n6708, \mem_REG.mem_2_22 , 
        n6707, \mem_REG.mem_2_21 , n6706, \mem_REG.mem_2_20 , n6705, 
        \mem_REG.mem_2_19 , n6704, \mem_REG.mem_2_18 , n6703, \mem_REG.mem_2_17 , 
        n6702, \mem_REG.mem_2_16 , n6701, \mem_REG.mem_2_15 , n6700, 
        \mem_REG.mem_2_14 , n6699, n6698, \mem_REG.mem_2_12 , n6697, 
        n6696, \mem_REG.mem_2_10 , n6695, n6694, n6693, \mem_REG.mem_2_7 , 
        n6692, \mem_REG.mem_2_6 , n6691, \mem_REG.mem_2_5 , n6690, 
        \mem_REG.mem_2_4 , n6689, \mem_REG.mem_2_3 , n6688, n6687, 
        \mem_REG.mem_2_1 , n6686, \mem_REG.mem_2_0 , n6685, \mem_REG.mem_1_31 , 
        n6684, \mem_REG.mem_1_30 , n6683, n6682, n6681, \mem_REG.mem_1_27 , 
        n6680, \mem_REG.mem_1_26 , n6679, n6678, n6677, \mem_REG.mem_1_23 , 
        n6676, \mem_REG.mem_1_22 , n6675, \mem_REG.mem_1_21 , n6674, 
        \mem_REG.mem_1_20 , n6673, \mem_REG.mem_1_19 , n6672, \mem_REG.mem_1_18 , 
        n6671, \mem_REG.mem_1_17 , n6670, \mem_REG.mem_1_16 , n6669, 
        \mem_REG.mem_1_15 , n6668, \mem_REG.mem_1_14 , n6667, n6666, 
        \mem_REG.mem_1_12 , n6665, n6664, \mem_REG.mem_1_10 , n6663, 
        n6662, n6661, \mem_REG.mem_1_7 , n6660, \mem_REG.mem_1_6 , 
        n6659, \mem_REG.mem_1_5 , n6658, \mem_REG.mem_1_4 , n6657, 
        \mem_REG.mem_1_3 , n6656, n6655, \mem_REG.mem_1_1 , n6654, 
        \mem_REG.mem_1_0 , n6653, \mem_REG.mem_0_31 , n6652, \mem_REG.mem_0_30 , 
        n6651, n6650, n6649, \mem_REG.mem_0_27 , n6648, \mem_REG.mem_0_26 , 
        n6647, n6646, n6645, \mem_REG.mem_0_23 , n6644, \mem_REG.mem_0_22 , 
        n6643, \mem_REG.mem_0_21 , n6642, \mem_REG.mem_0_20 , n6641, 
        \mem_REG.mem_0_19 , n6640, \mem_REG.mem_0_18 , n6639, \mem_REG.mem_0_17 , 
        n6638, \mem_REG.mem_0_16 , n6637, \mem_REG.mem_0_15 , n6636, 
        \mem_REG.mem_0_14 , n6635, n6634, \mem_REG.mem_0_12 , n6633, 
        n6632, \mem_REG.mem_0_10 , n6631, n6630, n6629, \mem_REG.mem_0_7 , 
        n6628, \mem_REG.mem_0_6 , n6627, \mem_REG.mem_0_5 , n6626, 
        \mem_REG.mem_0_4 , n6625, \mem_REG.mem_0_3 , n6624, n6623, 
        \mem_REG.mem_0_1 , n6622, \mem_REG.mem_0_0 , n15619, n9, n14509, 
        n14605, n7, n14608, n14905, n15589, n14512, n15577, n15559;
    wire [3:0]rd_addr_p1cmp_r;   // src/fifo_sc_32_lut_gen.v(125[48:63])
    
<<<<<<< Updated upstream
    FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_2 lscc_fifo_inst (.rd_fifo_en_w(rd_fifo_en_w), 
            .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r[7] ), .SLM_CLK_c(SLM_CLK_c), 
            .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r[6] ), .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r[5] ), 
            .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r[0] ), .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r[4] ), 
            .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r[3] ), .rd_addr_r({rd_addr_r}), 
            .reset_all_w(reset_all_w), .n8(n8), .wr_addr_r({wr_addr_r}), 
            .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r[2] ), .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r[1] ), 
            .GND_net(GND_net), .\rd_addr_p1_w[2] (\rd_addr_p1_w[2] ), .n14025(n14025), 
            .n6127(n6127), .VCC_net(VCC_net), .\fifo_temp_output[1] (\fifo_temp_output[1] ), 
            .n10430(n10430), .is_tx_fifo_full_flag(is_tx_fifo_full_flag), 
            .n6088(n6088), .\fifo_temp_output[0] (\fifo_temp_output[0] ), 
            .\wr_addr_p1_w[2] (\wr_addr_p1_w[2] ), .n1(n1), .n10226(n10226), 
            .n5989(n5989), .n5311(n5311), .\fifo_temp_output[4] (\fifo_temp_output[4] ), 
            .n5314(n5314), .\fifo_temp_output[5] (\fifo_temp_output[5] ), 
            .rx_buf_byte({rx_buf_byte}), .n5868(n5868), .n4882(n4882), 
            .\fifo_temp_output[2] (\fifo_temp_output[2] ), .n4887(n4887), 
            .\fifo_temp_output[3] (\fifo_temp_output[3] ), .n5536(n5536), 
            .\fifo_temp_output[6] (\fifo_temp_output[6] ), .n5539(n5539), 
            .\fifo_temp_output[7] (\fifo_temp_output[7] ), .n10786(n10786), 
            .is_fifo_empty_flag(is_fifo_empty_flag), .n4919(n4919), .n4922(n4922), 
            .fifo_write_cmd(fifo_write_cmd), .wr_fifo_en_w(wr_fifo_en_w), 
            .n4878(n4878), .rd_fifo_en_prev_r(rd_fifo_en_prev_r), .fifo_read_cmd(fifo_read_cmd)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_quad_word_mod.v(20[37:380])
>>>>>>> master
    
endmodule
//
// Verilog Description of module FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_3
//

module FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_3 (rd_addr_r, 
            SLM_CLK_c, reset_all_w, \mem_LUT.data_raw_r[0] , wr_addr_r, 
            fifo_write_cmd, is_tx_fifo_full_flag, wr_fifo_en_w, GND_net, 
            n2704, \wr_addr_p1_w[2] , n1, n10381, \mem_LUT.data_raw_r[7] , 
            \mem_LUT.data_raw_r[6] , \mem_LUT.data_raw_r[5] , \mem_LUT.data_raw_r[4] , 
            \mem_LUT.data_raw_r[3] , \mem_LUT.data_raw_r[2] , \mem_LUT.data_raw_r[1] , 
            rx_buf_byte, n5734, \fifo_temp_output[1] , n10640, VCC_net, 
            n5738, \fifo_temp_output[2] , n5633, rd_fifo_en_prev_r, 
            fifo_read_cmd, is_fifo_empty_flag, empty_o_N_1333, n11046, 
            n5741, \fifo_temp_output[3] , n5745, \fifo_temp_output[4] , 
            n5748, \fifo_temp_output[5] , n5812, \fifo_temp_output[0] , 
            n5755, \fifo_temp_output[6] , n5761, \fifo_temp_output[7] , 
            n5769, n5610, n5614, \rd_addr_p1_w[2] , n11863) /* synthesis syn_module_defined=1 */ ;
    output [2:0]rd_addr_r;
    input SLM_CLK_c;
    input reset_all_w;
    output \mem_LUT.data_raw_r[0] ;
    output [2:0]wr_addr_r;
    input fifo_write_cmd;
    output is_tx_fifo_full_flag;
    output wr_fifo_en_w;
    input GND_net;
    input n2704;
    output \wr_addr_p1_w[2] ;
    output n1;
    output n10381;
    output \mem_LUT.data_raw_r[7] ;
    output \mem_LUT.data_raw_r[6] ;
    output \mem_LUT.data_raw_r[5] ;
    output \mem_LUT.data_raw_r[4] ;
    output \mem_LUT.data_raw_r[3] ;
    output \mem_LUT.data_raw_r[2] ;
    output \mem_LUT.data_raw_r[1] ;
    input [7:0]rx_buf_byte;
    input n5734;
    output \fifo_temp_output[1] ;
    input n10640;
    input VCC_net;
    input n5738;
    output \fifo_temp_output[2] ;
    input n5633;
    output rd_fifo_en_prev_r;
    input fifo_read_cmd;
    output is_fifo_empty_flag;
    input empty_o_N_1333;
    input n11046;
    input n5741;
    output \fifo_temp_output[3] ;
    input n5745;
    output \fifo_temp_output[4] ;
    input n5748;
    output \fifo_temp_output[5] ;
    input n5812;
    output \fifo_temp_output[0] ;
    input n5755;
    output \fifo_temp_output[6] ;
    input n5761;
    output \fifo_temp_output[7] ;
    input n5769;
    input n5610;
    input n5614;
    output \rd_addr_p1_w[2] ;
    output n11863;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [2:0]n12;
    
    wire n11607, \mem_LUT.mem_1_1 , \mem_LUT.mem_0_1 ;
    wire [31:0]\mem_LUT.data_raw_r_31__N_1268 ;
    
    wire rd_fifo_en_w;
    wire [2:0]n12_adj_1365;
    
    wire \mem_LUT.mem_2_0 , \mem_LUT.mem_3_0 , n11613, n2, n11625, 
        \mem_LUT.mem_1_7 , \mem_LUT.mem_0_7 , \mem_LUT.mem_2_2 , \mem_LUT.mem_3_2 , 
        n11679, \mem_LUT.mem_1_2 , \mem_LUT.mem_0_2 , \mem_LUT.mem_2_3 , 
        \mem_LUT.mem_3_3 , n11673, \mem_LUT.mem_1_3 , \mem_LUT.mem_0_3 , 
        \mem_LUT.mem_2_1 , \mem_LUT.mem_3_1 , \mem_LUT.mem_1_0 , \mem_LUT.mem_0_0 , 
        \mem_LUT.mem_2_7 , \mem_LUT.mem_3_7 , \mem_LUT.mem_2_4 , \mem_LUT.mem_3_4 , 
        n11661, \mem_LUT.mem_1_4 , \mem_LUT.mem_0_4 , n3, n5806, \mem_LUT.mem_3_6 , 
        n5805, \mem_LUT.mem_3_5 , n5804, n5802, n5801, n5800, n5799, 
        n5797, \mem_LUT.mem_2_5 , n11655, \mem_LUT.mem_1_5 , \mem_LUT.mem_0_5 , 
        n4, n5796, \mem_LUT.mem_2_6 , n5795, n5794, n5793, n5792, 
        n5791, n5790, n5789, n5788, n5765, \mem_LUT.mem_1_6 , n5787, 
        n5786, n5785, n5784, n5783, n5782, n5779, n5778, n5777, 
        \mem_LUT.mem_0_6 , n5776, n5775, n5774, n5773, n5772, n5771, 
        n11637;
    
    SB_DFFSR rd_addr_r__i0 (.Q(rd_addr_r[0]), .C(SLM_CLK_c), .D(n12[0]), 
            .R(reset_all_w));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 n11607_bdd_4_lut (.I0(n11607), .I1(\mem_LUT.mem_1_1 ), .I2(\mem_LUT.mem_0_1 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1268 [1]));
    defparam n11607_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \mem_LUT.data_raw_r__i1  (.Q(\mem_LUT.data_raw_r[0] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1268 [0]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFSR wr_addr_r__i0 (.Q(wr_addr_r[0]), .C(SLM_CLK_c), .D(n12_adj_1365[0]), 
            .R(reset_all_w));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 wr_en_i_I_0_2_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(GND_net), .I3(GND_net), .O(wr_fifo_en_w));   // src/fifo_quad_word_mod.v(103[21:60])
    defparam wr_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1843_2_lut (.I0(wr_addr_r[0]), .I1(n2704), .I2(GND_net), 
            .I3(GND_net), .O(n12_adj_1365[0]));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1843_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10037 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_0 ), 
            .I2(\mem_LUT.mem_3_0 ), .I3(rd_addr_r[1]), .O(n11613));
    defparam rd_addr_r_0__bdd_4_lut_10037.LUT_INIT = 16'he4aa;
    SB_LUT4 i1619_3_lut (.I0(wr_addr_r[2]), .I1(wr_addr_r[1]), .I2(wr_addr_r[0]), 
            .I3(GND_net), .O(\wr_addr_p1_w[2] ));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam i1619_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1_4_lut (.I0(n1), .I1(\wr_addr_p1_w[2] ), .I2(n2), .I3(rd_addr_r[2]), 
            .O(n10381));
    defparam i1_4_lut.LUT_INIT = 16'h0208;
    SB_LUT4 wr_addr_r_1__I_0_i1_2_lut (.I0(wr_addr_r[0]), .I1(rd_addr_r[0]), 
            .I2(GND_net), .I3(GND_net), .O(n1));   // src/fifo_quad_word_mod.v(115[26:58])
    defparam wr_addr_r_1__I_0_i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n11625_bdd_4_lut (.I0(n11625), .I1(\mem_LUT.mem_1_7 ), .I2(\mem_LUT.mem_0_7 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1268 [7]));
    defparam n11625_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_2 ), 
            .I2(\mem_LUT.mem_3_2 ), .I3(rd_addr_r[1]), .O(n11679));
    defparam rd_addr_r_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n11679_bdd_4_lut (.I0(n11679), .I1(\mem_LUT.mem_1_2 ), .I2(\mem_LUT.mem_0_2 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1268 [2]));
    defparam n11679_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \mem_LUT.data_raw_r__i8  (.Q(\mem_LUT.data_raw_r[7] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1268 [7]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i7  (.Q(\mem_LUT.data_raw_r[6] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1268 [6]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i6  (.Q(\mem_LUT.data_raw_r[5] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1268 [5]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i5  (.Q(\mem_LUT.data_raw_r[4] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1268 [4]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i4  (.Q(\mem_LUT.data_raw_r[3] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1268 [3]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i3  (.Q(\mem_LUT.data_raw_r[2] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1268 [2]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i2  (.Q(\mem_LUT.data_raw_r[1] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1268 [1]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10081 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_3 ), 
            .I2(\mem_LUT.mem_3_3 ), .I3(rd_addr_r[1]), .O(n11673));
    defparam rd_addr_r_0__bdd_4_lut_10081.LUT_INIT = 16'he4aa;
    SB_LUT4 n11673_bdd_4_lut (.I0(n11673), .I1(\mem_LUT.mem_1_3 ), .I2(\mem_LUT.mem_0_3 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1268 [3]));
    defparam n11673_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10028 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_1 ), 
            .I2(\mem_LUT.mem_3_1 ), .I3(rd_addr_r[1]), .O(n11607));
    defparam rd_addr_r_0__bdd_4_lut_10028.LUT_INIT = 16'he4aa;
    SB_LUT4 n11613_bdd_4_lut (.I0(n11613), .I1(\mem_LUT.mem_1_0 ), .I2(\mem_LUT.mem_0_0 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1268 [0]));
    defparam n11613_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10047 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_7 ), 
            .I2(\mem_LUT.mem_3_7 ), .I3(rd_addr_r[1]), .O(n11625));
    defparam rd_addr_r_0__bdd_4_lut_10047.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10076 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_4 ), 
            .I2(\mem_LUT.mem_3_4 ), .I3(rd_addr_r[1]), .O(n11661));
    defparam rd_addr_r_0__bdd_4_lut_10076.LUT_INIT = 16'he4aa;
    SB_LUT4 n11661_bdd_4_lut (.I0(n11661), .I1(\mem_LUT.mem_1_4 ), .I2(\mem_LUT.mem_0_4 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1268 [4]));
    defparam n11661_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4347_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_3_7 ), .O(n5806));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4347_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4346_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_3_6 ), .O(n5805));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4346_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4345_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_3_5 ), .O(n5804));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4345_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF \mem_LUT.data_buff_r__i1  (.Q(\fifo_temp_output[1] ), .C(SLM_CLK_c), 
           .D(n5734));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 i4343_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_3_4 ), .O(n5802));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4343_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE full_r_84 (.Q(is_tx_fifo_full_flag), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n10640));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 i4342_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_3_3 ), .O(n5801));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4342_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_p1_w_1__I_0_i2_2_lut_3_lut (.I0(wr_addr_r[1]), .I1(wr_addr_r[0]), 
            .I2(rd_addr_r[1]), .I3(GND_net), .O(n2));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam wr_addr_p1_w_1__I_0_i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4341_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_3_2 ), .O(n5800));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4341_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4340_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_3_1 ), .O(n5799));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4340_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4338_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_3_0 ), .O(n5797));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4338_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10066 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_5 ), 
            .I2(\mem_LUT.mem_3_5 ), .I3(rd_addr_r[1]), .O(n11655));
    defparam rd_addr_r_0__bdd_4_lut_10066.LUT_INIT = 16'he4aa;
    SB_LUT4 n11655_bdd_4_lut (.I0(n11655), .I1(\mem_LUT.mem_1_5 ), .I2(\mem_LUT.mem_0_5 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1268 [5]));
    defparam n11655_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i3_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(GND_net), .O(n3));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i3_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF \mem_LUT.data_buff_r__i2  (.Q(\fifo_temp_output[2] ), .C(SLM_CLK_c), 
           .D(n5738));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 EnabledDecoder_2_i4_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(GND_net), .O(n4));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i4_2_lut_3_lut.LUT_INIT = 16'h0202;
<<<<<<< HEAD
    SB_LUT4 i4337_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_2_7 ), .O(n5796));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4337_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4336_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_2_6 ), .O(n5795));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4336_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4335_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_2_5 ), .O(n5794));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4335_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF rd_fifo_en_prev_r_86 (.Q(rd_fifo_en_prev_r), .C(SLM_CLK_c), .D(n5633));   // src/fifo_quad_word_mod.v(353[29] 363[32])
    SB_LUT4 i4334_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_2_4 ), .O(n5793));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4334_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4333_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_2_3 ), .O(n5792));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4333_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_en_i_I_0_2_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(GND_net), .I3(GND_net), .O(rd_fifo_en_w));   // src/fifo_quad_word_mod.v(62[29:51])
    defparam rd_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1846_2_lut (.I0(rd_addr_r[0]), .I1(empty_o_N_1333), .I2(GND_net), 
            .I3(GND_net), .O(n12[0]));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1846_2_lut.LUT_INIT = 16'h6666;
    SB_DFF empty_r_85 (.Q(is_fifo_empty_flag), .C(SLM_CLK_c), .D(n11046));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 i4332_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_2_2 ), .O(n5791));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4332_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4331_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_2_1 ), .O(n5790));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4331_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4330_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_2_0 ), .O(n5789));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4330_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF \mem_LUT.data_buff_r__i3  (.Q(\fifo_temp_output[3] ), .C(SLM_CLK_c), 
           .D(n5741));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i4  (.Q(\fifo_temp_output[4] ), .C(SLM_CLK_c), 
           .D(n5745));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i5  (.Q(\fifo_temp_output[5] ), .C(SLM_CLK_c), 
           .D(n5748));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE \mem_LUT.data_buff_r__i0  (.Q(\fifo_temp_output[0] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n5812));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i6  (.Q(\fifo_temp_output[6] ), .C(SLM_CLK_c), 
           .D(n5755));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 i4329_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_1_7 ), .O(n5788));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4329_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF \mem_LUT.data_buff_r__i7  (.Q(\fifo_temp_output[7] ), .C(SLM_CLK_c), 
           .D(n5761));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF i347_348 (.Q(\mem_LUT.mem_3_7 ), .C(SLM_CLK_c), .D(n5806));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i344_345 (.Q(\mem_LUT.mem_3_6 ), .C(SLM_CLK_c), .D(n5805));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i341_342 (.Q(\mem_LUT.mem_3_5 ), .C(SLM_CLK_c), .D(n5804));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF wr_addr_r__i1 (.Q(wr_addr_r[1]), .C(SLM_CLK_c), .D(n5765));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF i338_339 (.Q(\mem_LUT.mem_3_4 ), .C(SLM_CLK_c), .D(n5802));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i335_336 (.Q(\mem_LUT.mem_3_3 ), .C(SLM_CLK_c), .D(n5801));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i332_333 (.Q(\mem_LUT.mem_3_2 ), .C(SLM_CLK_c), .D(n5800));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i329_330 (.Q(\mem_LUT.mem_3_1 ), .C(SLM_CLK_c), .D(n5799));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF wr_addr_r__i2 (.Q(wr_addr_r[2]), .C(SLM_CLK_c), .D(n5769));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF i326_327 (.Q(\mem_LUT.mem_3_0 ), .C(SLM_CLK_c), .D(n5797));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i251_252 (.Q(\mem_LUT.mem_2_7 ), .C(SLM_CLK_c), .D(n5796));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i248_249 (.Q(\mem_LUT.mem_2_6 ), .C(SLM_CLK_c), .D(n5795));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i245_246 (.Q(\mem_LUT.mem_2_5 ), .C(SLM_CLK_c), .D(n5794));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i242_243 (.Q(\mem_LUT.mem_2_4 ), .C(SLM_CLK_c), .D(n5793));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i239_240 (.Q(\mem_LUT.mem_2_3 ), .C(SLM_CLK_c), .D(n5792));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i236_237 (.Q(\mem_LUT.mem_2_2 ), .C(SLM_CLK_c), .D(n5791));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i233_234 (.Q(\mem_LUT.mem_2_1 ), .C(SLM_CLK_c), .D(n5790));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i230_231 (.Q(\mem_LUT.mem_2_0 ), .C(SLM_CLK_c), .D(n5789));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i155_156 (.Q(\mem_LUT.mem_1_7 ), .C(SLM_CLK_c), .D(n5788));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 i4328_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_1_6 ), .O(n5787));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4328_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i152_153 (.Q(\mem_LUT.mem_1_6 ), .C(SLM_CLK_c), .D(n5787));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i149_150 (.Q(\mem_LUT.mem_1_5 ), .C(SLM_CLK_c), .D(n5786));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i146_147 (.Q(\mem_LUT.mem_1_4 ), .C(SLM_CLK_c), .D(n5785));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i143_144 (.Q(\mem_LUT.mem_1_3 ), .C(SLM_CLK_c), .D(n5784));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i140_141 (.Q(\mem_LUT.mem_1_2 ), .C(SLM_CLK_c), .D(n5783));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i137_138 (.Q(\mem_LUT.mem_1_1 ), .C(SLM_CLK_c), .D(n5782));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF rd_addr_r__i1 (.Q(rd_addr_r[1]), .C(SLM_CLK_c), .D(n5610));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF rd_addr_r__i2 (.Q(rd_addr_r[2]), .C(SLM_CLK_c), .D(n5614));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF i134_135 (.Q(\mem_LUT.mem_1_0 ), .C(SLM_CLK_c), .D(n5779));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i59_60 (.Q(\mem_LUT.mem_0_7 ), .C(SLM_CLK_c), .D(n5778));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i56_57 (.Q(\mem_LUT.mem_0_6 ), .C(SLM_CLK_c), .D(n5777));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i53_54 (.Q(\mem_LUT.mem_0_5 ), .C(SLM_CLK_c), .D(n5776));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i50_51 (.Q(\mem_LUT.mem_0_4 ), .C(SLM_CLK_c), .D(n5775));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 i4327_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_1_5 ), .O(n5786));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4327_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i47_48 (.Q(\mem_LUT.mem_0_3 ), .C(SLM_CLK_c), .D(n5774));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i44_45 (.Q(\mem_LUT.mem_0_2 ), .C(SLM_CLK_c), .D(n5773));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i41_42 (.Q(\mem_LUT.mem_0_1 ), .C(SLM_CLK_c), .D(n5772));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i38_39 (.Q(\mem_LUT.mem_0_0 ), .C(SLM_CLK_c), .D(n5771));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 i4326_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_1_4 ), .O(n5785));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4326_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4325_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_1_3 ), .O(n5784));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4325_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4324_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_1_2 ), .O(n5783));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4324_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4323_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_1_1 ), .O(n5782));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4323_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4320_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_1_0 ), .O(n5779));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4320_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4319_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_0_7 ), .O(n5778));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4319_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4318_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_0_6 ), .O(n5777));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4318_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4317_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_0_5 ), .O(n5776));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4317_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4306_4_lut_4_lut_4_lut (.I0(wr_addr_r[1]), .I1(wr_addr_r[0]), 
            .I2(n2704), .I3(reset_all_w), .O(n5765));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam i4306_4_lut_4_lut_4_lut.LUT_INIT = 16'h006a;
    SB_LUT4 i4316_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_0_4 ), .O(n5775));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4316_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10061 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_6 ), 
            .I2(\mem_LUT.mem_3_6 ), .I3(rd_addr_r[1]), .O(n11637));
    defparam rd_addr_r_0__bdd_4_lut_10061.LUT_INIT = 16'he4aa;
    SB_LUT4 i4315_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_0_3 ), .O(n5774));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4315_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4314_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_0_2 ), .O(n5773));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4314_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4313_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_0_1 ), .O(n5772));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4313_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4312_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_0_0 ), .O(n5771));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4312_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11637_bdd_4_lut (.I0(n11637), .I1(\mem_LUT.mem_1_6 ), .I2(\mem_LUT.mem_0_6 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1268 [6]));
    defparam n11637_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1641_3_lut (.I0(rd_addr_r[2]), .I1(rd_addr_r[1]), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(\rd_addr_p1_w[2] ));   // src/fifo_quad_word_mod.v(71[47:65])
    defparam i1641_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1634_rep_162_2_lut (.I0(rd_addr_r[1]), .I1(rd_addr_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n11863));   // src/fifo_quad_word_mod.v(71[47:65])
    defparam i1634_rep_162_2_lut.LUT_INIT = 16'h6666;
=======
    
endmodule
//
// Verilog Description of module spi
//

module spi (\tx_data_byte[3] , n2086, GND_net, \tx_data_byte[4] , SEN_c_1, 
            SLM_CLK_c, \tx_data_byte[5] , SOUT_c, n4312, \rx_shift_reg[0] , 
            \tx_data_byte[6] , n4319, SDAT_c_15, \tx_data_byte[7] , 
            tx_addr_byte, VCC_net, n10428, \tx_shift_reg[0] , n6060, 
            rx_buf_byte, n6059, n6058, n6057, n6056, n6055, n6054, 
            spi_rx_byte_ready, SCK_c_0, spi_start_transfer_r, n4897, 
            n4888, \rx_shift_reg[1] , n4883, \rx_shift_reg[2] , n4877, 
            \rx_shift_reg[3] , n4869, \rx_shift_reg[4] , n4838, \rx_shift_reg[5] , 
            multi_byte_spi_trans_flag_r, n4836, \rx_shift_reg[6] , n4834, 
            \rx_shift_reg[7] , \tx_data_byte[2] , \tx_data_byte[1] , n3495) /* synthesis syn_module_defined=1 */ ;
    input \tx_data_byte[3] ;
    output n2086;
    input GND_net;
    input \tx_data_byte[4] ;
    output SEN_c_1;
    input SLM_CLK_c;
    input \tx_data_byte[5] ;
    input SOUT_c;
    output n4312;
    output \rx_shift_reg[0] ;
    input \tx_data_byte[6] ;
    output n4319;
    output SDAT_c_15;
    input \tx_data_byte[7] ;
    input [7:0]tx_addr_byte;
    input VCC_net;
    input n10428;
    output \tx_shift_reg[0] ;
    input n6060;
    output [7:0]rx_buf_byte;
    input n6059;
    input n6058;
    input n6057;
    input n6056;
    input n6055;
    input n6054;
    output spi_rx_byte_ready;
    output SCK_c_0;
    input spi_start_transfer_r;
    input n4897;
    input n4888;
    output \rx_shift_reg[1] ;
    input n4883;
    output \rx_shift_reg[2] ;
    input n4877;
    output \rx_shift_reg[3] ;
    input n4869;
    output \rx_shift_reg[4] ;
    input n4838;
    output \rx_shift_reg[5] ;
    input multi_byte_spi_trans_flag_r;
    input n4836;
    output \rx_shift_reg[6] ;
    input n4834;
    output \rx_shift_reg[7] ;
    input \tx_data_byte[2] ;
    input \tx_data_byte[1] ;
    output n3495;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [15:0]tx_shift_reg;   // src/spi.v(70[12:24])
    wire [15:0]n2087;
    
    wire n7109;
    wire [3:0]state;   // src/spi.v(71[11:16])
    
    wire n12080;
    wire [9:0]counter;   // src/spi.v(69[11:18])
    
    wire n12081;
    wire [2:0]n970;
    wire [3:0]state_3__N_938;
    
    wire n10827, n24, n12108;
    wire [9:0]n45;
    
    wire n4380, n4694, n10203, n10204, n10202, n10201, n10200, 
        n10199, n10198, n10197, n10196;
    wire [7:0]n315;
    wire [7:0]multi_byte_counter;   // src/spi.v(68[11:29])
    wire [7:0]n2142;
    
    wire n10171, n10170, n10169, n10168, n10167, n10166, n10165, 
        n4, n37, n2, n4_adj_2, n51_adj_3, n12072, n3748, n12073, 
        n14, n19, n12052, n12057, n34, n37_adj_4, n10851, n4236, 
        n19_adj_5, n10778, n7, n4358, n10828, n10792, n10826, 
        n4_adj_6, n4629, n4541, n4672, n10, n14_adj_7, n34_adj_8, 
        n10_adj_9, n14_adj_10, n12101, n7_adj_11, n3, n3_adj_12, 
        n21, n10941, n22, n3_adj_13, n4519, n12112, n7_adj_14, 
        n12104;
    
    SB_LUT4 mux_981_i4_3_lut (.I0(\tx_data_byte[3] ), .I1(tx_shift_reg[2]), 
            .I2(n2086), .I3(GND_net), .O(n2087[3]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i5_3_lut (.I0(\tx_data_byte[4] ), .I1(tx_shift_reg[3]), 
            .I2(n2086), .I3(GND_net), .O(n2087[4]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10320_4_lut (.I0(n7109), .I1(state[1]), .I2(state[0]), .I3(state[2]), 
            .O(n12080));   // src/spi.v(88[9] 219[16])
    defparam i10320_4_lut.LUT_INIT = 16'hc08c;
    SB_LUT4 i1_4_lut (.I0(counter[4]), .I1(n12080), .I2(n12081), .I3(state[3]), 
            .O(n970[0]));   // src/spi.v(76[8] 221[4])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_DFF byte_recv_92_i2 (.Q(SEN_c_1), .C(SLM_CLK_c), .D(n970[1]));   // src/spi.v(88[9] 219[16])
    SB_LUT4 mux_981_i6_3_lut (.I0(\tx_data_byte[5] ), .I1(tx_shift_reg[4]), 
            .I2(n2086), .I3(GND_net), .O(n2087[5]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE rx_shift_reg_i0 (.Q(\rx_shift_reg[0] ), .C(SLM_CLK_c), .E(n4312), 
            .D(SOUT_c));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i0 (.Q(state[0]), .C(SLM_CLK_c), .E(n10827), .D(state_3__N_938[0]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i1_2_lut_3_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(GND_net), .O(n24));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i10319_2_lut_3_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(GND_net), .O(n12108));
    defparam i10319_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFFESR counter_1189__i0 (.Q(counter[0]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[0]), .R(n4694));   // src/spi.v(183[28:41])
    SB_LUT4 mux_981_i7_3_lut (.I0(\tx_data_byte[6] ), .I1(tx_shift_reg[5]), 
            .I2(n2086), .I3(GND_net), .O(n2087[6]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE tx_shift_reg_i0_i15 (.Q(SDAT_c_15), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[15]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_981_i8_3_lut (.I0(\tx_data_byte[7] ), .I1(tx_shift_reg[6]), 
            .I2(n2086), .I3(GND_net), .O(n2087[7]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i9_3_lut (.I0(tx_addr_byte[0]), .I1(tx_shift_reg[7]), 
            .I2(n2086), .I3(GND_net), .O(n2087[8]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i10_3_lut (.I0(tx_addr_byte[1]), .I1(tx_shift_reg[8]), 
            .I2(n2086), .I3(GND_net), .O(n2087[9]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i11_3_lut (.I0(tx_addr_byte[2]), .I1(tx_shift_reg[9]), 
            .I2(n2086), .I3(GND_net), .O(n2087[10]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i12_3_lut (.I0(tx_addr_byte[3]), .I1(tx_shift_reg[10]), 
            .I2(n2086), .I3(GND_net), .O(n2087[11]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i13_3_lut (.I0(tx_addr_byte[4]), .I1(tx_shift_reg[11]), 
            .I2(n2086), .I3(GND_net), .O(n2087[12]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i14_3_lut (.I0(tx_addr_byte[5]), .I1(tx_shift_reg[12]), 
            .I2(n2086), .I3(GND_net), .O(n2087[13]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i15_3_lut (.I0(tx_addr_byte[6]), .I1(tx_shift_reg[13]), 
            .I2(n2086), .I3(GND_net), .O(n2087[14]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY counter_1189_add_4_10 (.CI(n10203), .I0(VCC_net), .I1(counter[8]), 
            .CO(n10204));
    SB_LUT4 counter_1189_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[7]), 
            .I3(n10202), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFE tx_shift_reg_i0_i0 (.Q(\tx_shift_reg[0] ), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n10428));   // src/spi.v(76[8] 221[4])
    SB_CARRY counter_1189_add_4_9 (.CI(n10202), .I0(VCC_net), .I1(counter[7]), 
            .CO(n10203));
    SB_DFF Rx_Recv_Byte_i1 (.Q(rx_buf_byte[1]), .C(SLM_CLK_c), .D(n6060));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i2 (.Q(rx_buf_byte[2]), .C(SLM_CLK_c), .D(n6059));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i3 (.Q(rx_buf_byte[3]), .C(SLM_CLK_c), .D(n6058));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i4 (.Q(rx_buf_byte[4]), .C(SLM_CLK_c), .D(n6057));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i5 (.Q(rx_buf_byte[5]), .C(SLM_CLK_c), .D(n6056));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i6 (.Q(rx_buf_byte[6]), .C(SLM_CLK_c), .D(n6055));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i7 (.Q(rx_buf_byte[7]), .C(SLM_CLK_c), .D(n6054));   // src/spi.v(76[8] 221[4])
    SB_LUT4 counter_1189_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[6]), 
            .I3(n10201), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_8 (.CI(n10201), .I0(VCC_net), .I1(counter[6]), 
            .CO(n10202));
    SB_LUT4 counter_1189_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[5]), 
            .I3(n10200), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_7 (.CI(n10200), .I0(VCC_net), .I1(counter[5]), 
            .CO(n10201));
    SB_LUT4 counter_1189_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[4]), 
            .I3(n10199), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_6 (.CI(n10199), .I0(VCC_net), .I1(counter[4]), 
            .CO(n10200));
    SB_LUT4 counter_1189_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[3]), 
            .I3(n10198), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_5 (.CI(n10198), .I0(VCC_net), .I1(counter[3]), 
            .CO(n10199));
    SB_LUT4 counter_1189_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[2]), 
            .I3(n10197), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_4 (.CI(n10197), .I0(VCC_net), .I1(counter[2]), 
            .CO(n10198));
    SB_LUT4 counter_1189_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[1]), 
            .I3(n10196), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_3 (.CI(n10196), .I0(VCC_net), .I1(counter[1]), 
            .CO(n10197));
    SB_LUT4 counter_1189_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n10196));
    SB_LUT4 add_995_9_lut (.I0(GND_net), .I1(multi_byte_counter[7]), .I2(n2142[5]), 
            .I3(n10171), .O(n315[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_995_8_lut (.I0(GND_net), .I1(multi_byte_counter[6]), .I2(n2142[5]), 
            .I3(n10170), .O(n315[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_8 (.CI(n10170), .I0(multi_byte_counter[6]), .I1(n2142[5]), 
            .CO(n10171));
    SB_LUT4 add_995_7_lut (.I0(GND_net), .I1(multi_byte_counter[5]), .I2(n2142[5]), 
            .I3(n10169), .O(n315[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_7 (.CI(n10169), .I0(multi_byte_counter[5]), .I1(n2142[5]), 
            .CO(n10170));
    SB_LUT4 add_995_6_lut (.I0(GND_net), .I1(multi_byte_counter[4]), .I2(n2142[5]), 
            .I3(n10168), .O(n315[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_6 (.CI(n10168), .I0(multi_byte_counter[4]), .I1(n2142[5]), 
            .CO(n10169));
    SB_LUT4 add_995_5_lut (.I0(GND_net), .I1(multi_byte_counter[3]), .I2(n2142[5]), 
            .I3(n10167), .O(n315[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_5 (.CI(n10167), .I0(multi_byte_counter[3]), .I1(n2142[5]), 
            .CO(n10168));
    SB_LUT4 add_995_4_lut (.I0(GND_net), .I1(multi_byte_counter[2]), .I2(n2142[5]), 
            .I3(n10166), .O(n315[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_4 (.CI(n10166), .I0(multi_byte_counter[2]), .I1(n2142[5]), 
            .CO(n10167));
    SB_LUT4 add_995_3_lut (.I0(GND_net), .I1(multi_byte_counter[1]), .I2(n2142[5]), 
            .I3(n10165), .O(n315[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_3 (.CI(n10165), .I0(multi_byte_counter[1]), .I1(n2142[5]), 
            .CO(n10166));
    SB_LUT4 add_995_2_lut (.I0(GND_net), .I1(multi_byte_counter[0]), .I2(n2142[5]), 
            .I3(GND_net), .O(n315[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_2 (.CI(GND_net), .I0(multi_byte_counter[0]), .I1(n2142[5]), 
            .CO(n10165));
    SB_DFFE tx_shift_reg_i0_i14 (.Q(tx_shift_reg[14]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[14]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i13 (.Q(tx_shift_reg[13]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[13]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i12 (.Q(tx_shift_reg[12]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[12]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i11 (.Q(tx_shift_reg[11]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[11]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i10 (.Q(tx_shift_reg[10]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[10]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i9 (.Q(tx_shift_reg[9]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[9]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i8 (.Q(tx_shift_reg[8]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[8]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i7 (.Q(tx_shift_reg[7]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[7]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i6 (.Q(tx_shift_reg[6]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[6]));   // src/spi.v(76[8] 221[4])
    SB_DFF byte_recv_92_i3 (.Q(spi_rx_byte_ready), .C(SLM_CLK_c), .D(n970[2]));   // src/spi.v(88[9] 219[16])
    SB_DFFE tx_shift_reg_i0_i5 (.Q(tx_shift_reg[5]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[5]));   // src/spi.v(76[8] 221[4])
    SB_DFF byte_recv_92_i1 (.Q(SCK_c_0), .C(SLM_CLK_c), .D(n970[0]));   // src/spi.v(88[9] 219[16])
    SB_DFFE tx_shift_reg_i0_i4 (.Q(tx_shift_reg[4]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[4]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i3 (.Q(tx_shift_reg[3]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[3]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i1_2_lut (.I0(state[3]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n4));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_3 (.I0(n37), .I1(state[0]), .I2(n2), .I3(n4_adj_2), 
            .O(n2086));
    defparam i1_4_lut_adj_3.LUT_INIT = 16'ha2a0;
    SB_LUT4 i1_2_lut_adj_4 (.I0(counter[4]), .I1(n51_adj_3), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // src/spi.v(183[28:41])
    defparam i1_2_lut_adj_4.LUT_INIT = 16'h4444;
    SB_LUT4 i10314_4_lut (.I0(spi_start_transfer_r), .I1(state[0]), .I2(n37), 
            .I3(state[3]), .O(n12072));   // src/spi.v(71[11:16])
    defparam i10314_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1_4_lut_adj_5 (.I0(n3748), .I1(n12072), .I2(n12073), .I3(state[1]), 
            .O(n4319));
    defparam i1_4_lut_adj_5.LUT_INIT = 16'h5044;
    SB_LUT4 mux_981_i16_3_lut (.I0(tx_addr_byte[7]), .I1(tx_shift_reg[14]), 
            .I2(n2086), .I3(GND_net), .O(n2087[15]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(state[3]), .I1(state[2]), .I2(state[0]), .I3(GND_net), 
            .O(n14));   // src/spi.v(88[9] 219[16])
    defparam i1_3_lut.LUT_INIT = 16'hcdcd;
    SB_LUT4 i10301_3_lut (.I0(state[0]), .I1(state[2]), .I2(n19), .I3(GND_net), 
            .O(n12052));
    defparam i10301_3_lut.LUT_INIT = 16'h4d4d;
    SB_LUT4 i10298_3_lut (.I0(state[3]), .I1(state[2]), .I2(state[0]), 
            .I3(GND_net), .O(n12057));
    defparam i10298_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF Rx_Recv_Byte_i0 (.Q(rx_buf_byte[0]), .C(SLM_CLK_c), .D(n4897));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i65_3_lut (.I0(n14), .I1(n12052), .I2(state[1]), .I3(GND_net), 
            .O(n34));
    defparam i65_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i66_4_lut (.I0(n12057), .I1(n2142[5]), .I2(state[1]), .I3(state[3]), 
            .O(n37_adj_4));
    defparam i66_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_4_lut_adj_6 (.I0(state[3]), .I1(n37_adj_4), .I2(n34), .I3(n10851), 
            .O(n4694));
    defparam i1_4_lut_adj_6.LUT_INIT = 16'h50dc;
    SB_LUT4 i10430_4_lut (.I0(state[3]), .I1(state[1]), .I2(n4236), .I3(n14), 
            .O(n4380));   // src/spi.v(88[9] 219[16])
    defparam i10430_4_lut.LUT_INIT = 16'h4c5f;
    SB_DFF rx_shift_reg_i1 (.Q(\rx_shift_reg[1] ), .C(SLM_CLK_c), .D(n4888));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i2 (.Q(tx_shift_reg[2]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[2]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i1 (.Q(tx_shift_reg[1]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[1]));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i2 (.Q(\rx_shift_reg[2] ), .C(SLM_CLK_c), .D(n4883));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i3 (.Q(state[3]), .C(SLM_CLK_c), .E(n19_adj_5), .D(state_3__N_938[3]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i2_3_lut (.I0(state[3]), .I1(n19), .I2(state[1]), .I3(GND_net), 
            .O(n10778));
    defparam i2_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i4_4_lut (.I0(n7), .I1(state[3]), .I2(spi_start_transfer_r), 
            .I3(state[0]), .O(n4358));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(state[1]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n7));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFFE state_i2 (.Q(state[2]), .C(SLM_CLK_c), .E(n10828), .D(state_3__N_938[2]));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i1 (.Q(state[1]), .C(SLM_CLK_c), .E(n10792), .D(state_3__N_938[1]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i1_4_lut_adj_7 (.I0(n4358), .I1(n10778), .I2(state[0]), .I3(state[2]), 
            .O(n10826));
    defparam i1_4_lut_adj_7.LUT_INIT = 16'h8aaa;
    SB_DFF rx_shift_reg_i3 (.Q(\rx_shift_reg[3] ), .C(SLM_CLK_c), .D(n4877));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i1_2_lut_adj_8 (.I0(n19), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_6));
    defparam i1_2_lut_adj_8.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_4_lut_adj_9 (.I0(state[3]), .I1(n10826), .I2(n7), .I3(n4_adj_6), 
            .O(n10827));
    defparam i1_4_lut_adj_9.LUT_INIT = 16'h4c44;
    SB_LUT4 i3_4_lut (.I0(counter[0]), .I1(counter[3]), .I2(counter[2]), 
            .I3(counter[1]), .O(n51_adj_3));   // src/spi.v(183[28:41])
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i9015_2_lut (.I0(state[0]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n10851));
    defparam i9015_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_10 (.I0(state[2]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n3748));   // src/spi.v(88[9] 219[16])
    defparam i1_2_lut_adj_10.LUT_INIT = 16'h2222;
    SB_LUT4 i10440_3_lut (.I0(counter[4]), .I1(n4629), .I2(n51_adj_3), 
            .I3(GND_net), .O(n4312));   // src/spi.v(88[9] 219[16])
    defparam i10440_3_lut.LUT_INIT = 16'h2020;
    SB_DFFESR counter_1189__i1 (.Q(counter[1]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[1]), .R(n4694));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1189__i2 (.Q(counter[2]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[2]), .R(n4694));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1189__i3 (.Q(counter[3]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[3]), .R(n4694));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1189__i4 (.Q(counter[4]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[4]), .R(n4694));   // src/spi.v(183[28:41])
    SB_DFF rx_shift_reg_i4 (.Q(\rx_shift_reg[4] ), .C(SLM_CLK_c), .D(n4869));   // src/spi.v(76[8] 221[4])
    SB_DFFESR counter_1189__i5 (.Q(counter[5]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[5]), .R(n4694));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1189__i9 (.Q(counter[9]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[9]), .R(n4694));   // src/spi.v(183[28:41])
    SB_DFFESS counter_1189__i8 (.Q(counter[8]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[8]), .S(n4694));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1189__i7 (.Q(counter[7]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[7]), .R(n4694));   // src/spi.v(183[28:41])
    SB_DFFESR multi_byte_counter_i1 (.Q(multi_byte_counter[1]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[1]), .R(n4672));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i2 (.Q(multi_byte_counter[2]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[2]), .R(n4672));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i3 (.Q(multi_byte_counter[3]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[3]), .R(n4672));   // src/spi.v(76[8] 221[4])
    SB_DFFESR counter_1189__i6 (.Q(counter[6]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[6]), .R(n4694));   // src/spi.v(183[28:41])
    SB_DFFESR multi_byte_counter_i4 (.Q(multi_byte_counter[4]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[4]), .R(n4672));   // src/spi.v(76[8] 221[4])
    SB_DFFESS multi_byte_counter_i5 (.Q(multi_byte_counter[5]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[5]), .S(n4672));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i2_2_lut_adj_11 (.I0(multi_byte_counter[2]), .I1(multi_byte_counter[4]), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // src/spi.v(208[21:52])
    defparam i2_2_lut_adj_11.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(multi_byte_counter[3]), .I1(multi_byte_counter[1]), 
            .I2(multi_byte_counter[5]), .I3(multi_byte_counter[7]), .O(n14_adj_7));   // src/spi.v(208[21:52])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(multi_byte_counter[0]), .I1(n14_adj_7), .I2(n10), 
            .I3(multi_byte_counter[6]), .O(n2142[5]));   // src/spi.v(208[21:52])
    defparam i7_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i2_3_lut_adj_12 (.I0(counter[2]), .I1(counter[1]), .I2(counter[3]), 
            .I3(GND_net), .O(n34_adj_8));   // src/spi.v(183[28:41])
    defparam i2_3_lut_adj_12.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_2_lut_adj_13 (.I0(counter[6]), .I1(counter[7]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_9));   // src/spi.v(141[21:41])
    defparam i2_2_lut_adj_13.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_14 (.I0(counter[4]), .I1(counter[5]), .I2(counter[9]), 
            .I3(n34_adj_8), .O(n14_adj_10));   // src/spi.v(141[21:41])
    defparam i6_4_lut_adj_14.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_15 (.I0(counter[0]), .I1(n14_adj_10), .I2(n10_adj_9), 
            .I3(counter[8]), .O(n19));   // src/spi.v(141[21:41])
    defparam i7_4_lut_adj_15.LUT_INIT = 16'hfffd;
    SB_LUT4 i10345_3_lut (.I0(n2142[5]), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n12101));   // src/spi.v(88[9] 219[16])
    defparam i10345_3_lut.LUT_INIT = 16'hc4c4;
    SB_LUT4 mux_344_Mux_1_i7_4_lut (.I0(state[0]), .I1(state[2]), .I2(n19), 
            .I3(state[1]), .O(n7_adj_11));   // src/spi.v(88[9] 219[16])
    defparam mux_344_Mux_1_i7_4_lut.LUT_INIT = 16'h02dd;
    SB_LUT4 mux_344_Mux_1_i15_4_lut (.I0(n7_adj_11), .I1(n12101), .I2(state[3]), 
            .I3(state[2]), .O(n970[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_344_Mux_1_i15_4_lut.LUT_INIT = 16'hfaca;
    SB_DFFESR multi_byte_counter_i0 (.Q(multi_byte_counter[0]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[0]), .R(n4672));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i6 (.Q(multi_byte_counter[6]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[6]), .R(n4672));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i5 (.Q(\rx_shift_reg[5] ), .C(SLM_CLK_c), .D(n4838));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_56_Mux_1_i3_3_lut_3_lut (.I0(multi_byte_spi_trans_flag_r), 
            .I1(state[0]), .I2(state[1]), .I3(GND_net), .O(n3));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_1_i3_3_lut_3_lut.LUT_INIT = 16'h3e3e;
    SB_LUT4 mux_56_Mux_0_i3_4_lut_4_lut (.I0(multi_byte_spi_trans_flag_r), 
            .I1(state[0]), .I2(state[1]), .I3(n19), .O(n3_adj_12));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_0_i3_4_lut_4_lut.LUT_INIT = 16'hc131;
    SB_DFFESS multi_byte_counter_i7 (.Q(multi_byte_counter[7]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[7]), .S(n4672));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i6 (.Q(\rx_shift_reg[6] ), .C(SLM_CLK_c), .D(n4836));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i43_4_lut_4_lut (.I0(state[3]), .I1(state[2]), .I2(state[1]), 
            .I3(state[0]), .O(n21));
    defparam i43_4_lut_4_lut.LUT_INIT = 16'hf01a;
    SB_LUT4 i3273_3_lut_4_lut (.I0(state[3]), .I1(state[2]), .I2(state[0]), 
            .I3(n3_adj_12), .O(state_3__N_938[0]));
    defparam i3273_3_lut_4_lut.LUT_INIT = 16'h1f0e;
    SB_DFF rx_shift_reg_i7 (.Q(\rx_shift_reg[7] ), .C(SLM_CLK_c), .D(n4834));   // src/spi.v(76[8] 221[4])
    SB_LUT4 counter_1189_add_4_11_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[9]), 
            .I3(n10204), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1189_add_4_10_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[8]), 
            .I3(n10203), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_981_i3_3_lut (.I0(\tx_data_byte[2] ), .I1(tx_shift_reg[1]), 
            .I2(n2086), .I3(GND_net), .O(n2087[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i2_3_lut (.I0(\tx_data_byte[1] ), .I1(\tx_shift_reg[0] ), 
            .I2(n2086), .I3(GND_net), .O(n2087[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[2]), .I1(n10778), .I2(n4358), .I3(state[0]), 
            .O(n10828));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hc0e0;
    SB_LUT4 i9104_3_lut_4_lut (.I0(state[0]), .I1(state[2]), .I2(spi_start_transfer_r), 
            .I3(state[1]), .O(n10941));
    defparam i9104_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_56_Mux_3_i15_4_lut (.I0(n12108), .I1(state[1]), .I2(state[3]), 
            .I3(n2142[5]), .O(state_3__N_938[3]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_3_i15_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i10427_4_lut (.I0(n22), .I1(n10941), .I2(n24), .I3(state[3]), 
            .O(n19_adj_5));
    defparam i10427_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i1_2_lut_adj_16 (.I0(n19), .I1(n21), .I2(GND_net), .I3(GND_net), 
            .O(n22));
    defparam i1_2_lut_adj_16.LUT_INIT = 16'h8888;
    SB_LUT4 i10306_2_lut_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(n7109), .O(n12081));   // src/spi.v(88[9] 219[16])
    defparam i10306_2_lut_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 mux_56_Mux_2_i15_4_lut (.I0(n3_adj_13), .I1(state[2]), .I2(state[3]), 
            .I3(state[0]), .O(state_3__N_938[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_2_i15_4_lut.LUT_INIT = 16'hc2ce;
    SB_LUT4 mux_56_Mux_2_i3_3_lut (.I0(multi_byte_spi_trans_flag_r), .I1(state[0]), 
            .I2(state[1]), .I3(GND_net), .O(n3_adj_13));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_2_i3_3_lut.LUT_INIT = 16'hc2c2;
    SB_LUT4 i1_2_lut_adj_17 (.I0(state[2]), .I1(n10778), .I2(GND_net), 
            .I3(GND_net), .O(n4519));
    defparam i1_2_lut_adj_17.LUT_INIT = 16'heeee;
    SB_LUT4 mux_56_Mux_1_i7_4_lut (.I0(n3), .I1(n12112), .I2(state[2]), 
            .I3(state[1]), .O(n7_adj_14));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_1_i7_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i2050_4_lut_4_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(state[3]), .O(n4629));   // src/spi.v(88[9] 219[16])
    defparam i2050_4_lut_4_lut_4_lut.LUT_INIT = 16'hfe75;
    SB_LUT4 i10352_2_lut (.I0(n19), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n12112));   // src/spi.v(88[9] 219[16])
    defparam i10352_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_4_lut (.I0(state[3]), .I1(n4519), .I2(n24), .I3(n4358), 
            .O(n10792));
    defparam i2_4_lut.LUT_INIT = 16'h4c00;
    SB_LUT4 i1_4_lut_adj_18 (.I0(state[1]), .I1(n4), .I2(n12104), .I3(state[0]), 
            .O(n4541));
    defparam i1_4_lut_adj_18.LUT_INIT = 16'ha088;
    SB_LUT4 i10290_3_lut (.I0(state[3]), .I1(state[2]), .I2(n19), .I3(GND_net), 
            .O(n12104));
    defparam i10290_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i3289_2_lut (.I0(n4541), .I1(state[3]), .I2(GND_net), .I3(GND_net), 
            .O(n4672));   // src/spi.v(76[8] 221[4])
    defparam i3289_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_4_lut (.I0(n2142[5]), .I1(state[0]), .I2(state[2]), 
            .I3(state[1]), .O(n4236));   // src/spi.v(88[9] 219[16])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[0]), .I1(state[2]), .I2(state[1]), 
            .I3(state[3]), .O(n2));   // src/spi.v(88[9] 219[16])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h00b0;
    SB_LUT4 i10326_2_lut_3_lut (.I0(counter[4]), .I1(n51_adj_3), .I2(state[3]), 
            .I3(GND_net), .O(n12073));   // src/spi.v(71[11:16])
    defparam i10326_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_3_lut_adj_19 (.I0(state[1]), .I1(state[3]), .I2(state[2]), 
            .I3(GND_net), .O(n4_adj_2));
    defparam i1_2_lut_3_lut_adj_19.LUT_INIT = 16'h0404;
    SB_LUT4 i2123_4_lut_4_lut (.I0(state[0]), .I1(state[2]), .I2(state[1]), 
            .I3(state[3]), .O(n3495));   // src/spi.v(88[9] 219[16])
    defparam i2123_4_lut_4_lut.LUT_INIT = 16'hfdfb;
    SB_LUT4 mux_344_Mux_2_i15_4_lut_4_lut (.I0(state[0]), .I1(state[1]), 
            .I2(state[2]), .I3(state[3]), .O(n970[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_344_Mux_2_i15_4_lut_4_lut.LUT_INIT = 16'h0420;
    SB_LUT4 mux_56_Mux_1_i15_3_lut_4_lut (.I0(state[0]), .I1(state[1]), 
            .I2(state[3]), .I3(n7_adj_14), .O(state_3__N_938[1]));
    defparam mux_56_Mux_1_i15_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i1_2_lut_4_lut_adj_20 (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(counter[3]), .O(n7109));   // src/spi.v(183[28:41])
    defparam i1_2_lut_4_lut_adj_20.LUT_INIT = 16'hfffe;
=======
    wire n3679, n3402;
    wire [3:0]n2775;
    
    wire n3400, n2, n4, n13687, n13688, n15499, n3398, n2057, 
        n13676, n13675, n12302, n13714, n13715, n15475, n4_adj_1365, 
        n14587, n12301, n6_adj_1366, n12968, n12990, \MISC.wr_w , 
        n13046, full_nxt_w_N_812, empty_nxt_w_N_823, n13700, n13699, 
        n14590, n4_adj_1367;
    wire [3:0]wr_addr_p1_r;   // src/fifo_sc_32_lut_gen.v(118[48:60])
    wire [2:0]wr_cmpaddr_p1_r;   // src/fifo_sc_32_lut_gen.v(122[54:69])
    
    wire n6_adj_1368, n12972, full_nxt_w_N_797, n12934;
    wire [3:0]rd_addr_nxt_w;   // src/fifo_sc_32_lut_gen.v(133[28:41])
    wire [31:0]sc32_fifo_data_out;   // src/top.v(613[12:30])
    
    wire n14737, n14740, n13132, n13133, n14731, n13130, n13129, 
        n13663, n13664, n15451, n13646, n13645;
    wire [3:0]wr_addr_nxt_w;   // src/fifo_sc_32_lut_gen.v(130[28:41])
    
    wire n13813, n13814, n15433, n13637, n13636, n13702, n13703, 
        n15409, n13622, n13621, n16201, n16204;
    wire [3:0]wr_addr_p1cmp_r_3__N_698;
    
    wire n16159, n16162, n13816, n13817, n15373, n13574, n13573, 
        n16063, n16066, n15283, n15286, n15259, n15262, n15985, 
        n15988, n15211, n15214, n15193, n14569, n15196, n14203, 
        n14204, n15925, n14192, n14191, n14185, n14186, n15919, 
        n14168, n14167, n14572, n15121, n15124, n15853, n15856, 
        n15835, n15838, n15811, n15814, n13456, n13457, n15079, 
        n13334, n13333, n15799, n15802, n3090, n3119;
    
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_13466  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_28 ), .I2(\mem_REG.mem_3_28 ), .I3(rd_addr_r[1]), 
            .O(n15781));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_13466 .LUT_INIT = 16'he4aa;
    SB_LUT4 n15781_bdd_4_lut (.I0(n15781), .I1(\mem_REG.mem_1_28 ), .I2(\mem_REG.mem_0_28 ), 
            .I3(rd_addr_r[1]), .O(n15784));
    defparam n15781_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_12582  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_13 ), .I2(\mem_REG.mem_3_13 ), .I3(rd_addr_r[1]), 
            .O(n14635));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_12582 .LUT_INIT = 16'he4aa;
    SB_DFFE \mem_REG.data_raw_r_i0_i1  (.Q(DEBUG_9_c_0), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[0]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_LUT4 n14635_bdd_4_lut (.I0(n14635), .I1(\mem_REG.mem_1_13 ), .I2(\mem_REG.mem_0_13 ), 
            .I3(rd_addr_r[1]), .O(n14638));
    defparam n14635_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_13451  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_28 ), .I2(\mem_REG.mem_7_28 ), .I3(rd_addr_r[1]), 
            .O(n15739));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_13451 .LUT_INIT = 16'he4aa;
    SB_LUT4 n15739_bdd_4_lut (.I0(n15739), .I1(\mem_REG.mem_5_28 ), .I2(\mem_REG.mem_4_28 ), 
            .I3(rd_addr_r[1]), .O(n15742));
    defparam n15739_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13566 (.I0(rd_addr_r[1]), .I1(n13801), 
            .I2(n13802), .I3(rd_addr_r[2]), .O(n15733));
    defparam rd_addr_r_1__bdd_4_lut_13566.LUT_INIT = 16'he4aa;
    SB_LUT4 n15733_bdd_4_lut (.I0(n15733), .I1(n13781), .I2(n13780), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[10]));
    defparam n15733_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13411 (.I0(rd_addr_r[1]), .I1(n13807), 
            .I2(n13808), .I3(rd_addr_r[2]), .O(n15727));
    defparam rd_addr_r_1__bdd_4_lut_13411.LUT_INIT = 16'he4aa;
    SB_LUT4 n15727_bdd_4_lut (.I0(n15727), .I1(n13784), .I2(n13783), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[27]));
    defparam n15727_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5403_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[31] ), 
            .I3(\mem_REG.mem_7_31 ), .O(n6877));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5403_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5402_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[30] ), 
            .I3(\mem_REG.mem_7_30 ), .O(n6876));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5402_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5401_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[29] ), 
            .I3(\mem_REG.mem_7_29 ), .O(n6875));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5401_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF \MISC.wr_flag_addr_r_i0  (.Q(\MISC.wr_flag_addr_r [0]), .C(SLM_CLK_c), 
           .D(wr_addr_r_3__N_690[0]));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_DFF \MISC.wr_flag_addr_p1_r_i0  (.Q(\MISC.wr_flag_addr_p1_r [0]), .C(SLM_CLK_c), 
           .D(wr_addr_p1_r_3__N_694[0]));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_LUT4 i5400_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[28] ), 
            .I3(\mem_REG.mem_7_28 ), .O(n6874));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5400_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF \MISC.rd_flag_addr_r_i0  (.Q(\MISC.rd_flag_addr_r [0]), .C(SLM_CLK_c), 
           .D(rd_addr_r_3__N_708[0]));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_LUT4 i5399_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[27] ), 
            .I3(\mem_REG.mem_7_27 ), .O(n6873));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5399_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5398_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[26] ), 
            .I3(\mem_REG.mem_7_26 ), .O(n6872));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5398_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5397_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[25] ), 
            .I3(\mem_REG.mem_7_25 ), .O(n6871));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5397_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF \MISC.rd_flag_addr_p1_r_i0  (.Q(\MISC.rd_flag_addr_p1_r [0]), .C(SLM_CLK_c), 
           .D(rd_addr_p1_r_3__N_712[0]));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_LUT4 i5396_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[24] ), 
            .I3(\mem_REG.mem_7_24 ), .O(n6870));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5396_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF \MISC.full_flag_r_143  (.Q(\MISC.full_flag_r ), .C(SLM_CLK_c), 
           .D(full_ext_r_N_794));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_DFF \MISC.empty_flag_r_144  (.Q(\MISC.empty_flag_r ), .C(SLM_CLK_c), 
           .D(empty_ext_r_N_796));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_LUT4 i5395_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[23] ), 
            .I3(\mem_REG.mem_7_23 ), .O(n6869));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5395_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFSS \MISC.AEmpty.almost_empty_ext_r_147  (.Q(sc32_fifo_almost_empty), 
            .C(SLM_CLK_c), .D(\MISC.AEmpty.almost_empty_nxt_w ), .S(reset_all));   // src/fifo_sc_32_lut_gen.v(403[33] 415[36])
    SB_LUT4 i5394_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[22] ), 
            .I3(\mem_REG.mem_7_22 ), .O(n6868));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5394_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5393_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[21] ), 
            .I3(\mem_REG.mem_7_21 ), .O(n6867));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5393_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5392_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[20] ), 
            .I3(\mem_REG.mem_7_20 ), .O(n6866));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5392_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5391_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[19] ), 
            .I3(\mem_REG.mem_7_19 ), .O(n6865));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5391_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5390_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[18] ), 
            .I3(\mem_REG.mem_7_18 ), .O(n6864));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5390_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5389_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[17] ), 
            .I3(\mem_REG.mem_7_17 ), .O(n6863));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5389_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5388_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[16] ), 
            .I3(\mem_REG.mem_7_16 ), .O(n6862));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5388_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12867 (.I0(rd_addr_r[1]), .I1(n13723), 
            .I2(n13724), .I3(rd_addr_r[2]), .O(n15001));
    defparam rd_addr_r_1__bdd_4_lut_12867.LUT_INIT = 16'he4aa;
    SB_LUT4 i5387_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[15] ), 
            .I3(\mem_REG.mem_7_15 ), .O(n6861));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5387_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5386_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[14] ), 
            .I3(\mem_REG.mem_7_14 ), .O(n6860));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5386_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5385_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[13] ), 
            .I3(\mem_REG.mem_7_13 ), .O(n6859));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5385_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5384_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[12] ), 
            .I3(\mem_REG.mem_7_12 ), .O(n6858));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5384_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15001_bdd_4_lut (.I0(n15001), .I1(n13430), .I2(n13429), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[19]));
    defparam n15001_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5383_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[11] ), 
            .I3(\mem_REG.mem_7_11 ), .O(n6857));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5383_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5382_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[10] ), 
            .I3(\mem_REG.mem_7_10 ), .O(n6856));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5382_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5381_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[9] ), 
            .I3(\mem_REG.mem_7_9 ), .O(n6855));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5381_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5380_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[8] ), 
            .I3(\mem_REG.mem_7_8 ), .O(n6854));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5380_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_13416  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_11 ), .I2(\mem_REG.mem_3_11 ), .I3(rd_addr_r[1]), 
            .O(n15703));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_13416 .LUT_INIT = 16'he4aa;
    SB_LUT4 i5379_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[7] ), 
            .I3(\mem_REG.mem_7_7 ), .O(n6853));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5379_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15703_bdd_4_lut (.I0(n15703), .I1(\mem_REG.mem_1_11 ), .I2(\mem_REG.mem_0_11 ), 
            .I3(rd_addr_r[1]), .O(n15706));
    defparam n15703_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_13386  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_1 ), .I2(\mem_REG.mem_7_1 ), .I3(rd_addr_r[1]), 
            .O(n15697));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_13386 .LUT_INIT = 16'he4aa;
    SB_LUT4 n15697_bdd_4_lut (.I0(n15697), .I1(\mem_REG.mem_5_1 ), .I2(\mem_REG.mem_4_1 ), 
            .I3(rd_addr_r[1]), .O(n15700));
    defparam n15697_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5378_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[6] ), 
            .I3(\mem_REG.mem_7_6 ), .O(n6852));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5378_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11567_3_lut (.I0(\mem_REG.mem_0_8 ), .I1(\mem_REG.mem_1_8 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13678));
    defparam i11567_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11568_3_lut (.I0(\mem_REG.mem_2_8 ), .I1(\mem_REG.mem_3_8 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13679));
    defparam i11568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5377_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[5] ), 
            .I3(\mem_REG.mem_7_5 ), .O(n6851));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5377_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11598_3_lut (.I0(\mem_REG.mem_6_8 ), .I1(\mem_REG.mem_7_8 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13709));
    defparam i11598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11597_3_lut (.I0(\mem_REG.mem_4_8 ), .I1(\mem_REG.mem_5_8 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13708));
    defparam i11597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5376_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[4] ), 
            .I3(\mem_REG.mem_7_4 ), .O(n6850));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5376_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5375_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[3] ), 
            .I3(\mem_REG.mem_7_3 ), .O(n6849));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5375_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12802 (.I0(rd_addr_r[1]), .I1(n13732), 
            .I2(n13733), .I3(rd_addr_r[2]), .O(n14983));
    defparam rd_addr_r_1__bdd_4_lut_12802.LUT_INIT = 16'he4aa;
    SB_LUT4 i5374_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[2] ), 
            .I3(\mem_REG.mem_7_2 ), .O(n6848));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5374_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5373_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[1] ), 
            .I3(\mem_REG.mem_7_1 ), .O(n6847));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5373_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14983_bdd_4_lut (.I0(n14983), .I1(n13151), .I2(n13150), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[18]));
    defparam n14983_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5372_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(DEBUG_5_c_0), 
            .I3(\mem_REG.mem_7_0 ), .O(n6846));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5372_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11609_3_lut (.I0(\mem_REG.mem_0_24 ), .I1(\mem_REG.mem_1_24 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13720));
    defparam i11609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11610_3_lut (.I0(\mem_REG.mem_2_24 ), .I1(\mem_REG.mem_3_24 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13721));
    defparam i11610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11616_3_lut (.I0(\mem_REG.mem_6_24 ), .I1(\mem_REG.mem_7_24 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13727));
    defparam i11616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11615_3_lut (.I0(\mem_REG.mem_4_24 ), .I1(\mem_REG.mem_5_24 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13726));
    defparam i11615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11633_3_lut (.I0(\mem_REG.mem_0_9 ), .I1(\mem_REG.mem_1_9 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13744));
    defparam i11633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11634_3_lut (.I0(\mem_REG.mem_2_9 ), .I1(\mem_REG.mem_3_9 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13745));
    defparam i11634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11694_3_lut (.I0(\mem_REG.mem_6_9 ), .I1(\mem_REG.mem_7_9 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13805));
    defparam i11694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11693_3_lut (.I0(\mem_REG.mem_4_9 ), .I1(\mem_REG.mem_5_9 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13804));
    defparam i11693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11216_3_lut (.I0(\mem_REG.mem_0_2 ), .I1(\mem_REG.mem_1_2 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13327));
    defparam i11216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11217_3_lut (.I0(\mem_REG.mem_2_2 ), .I1(\mem_REG.mem_3_2 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13328));
    defparam i11217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11220_3_lut (.I0(\mem_REG.mem_6_2 ), .I1(\mem_REG.mem_7_2 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13331));
    defparam i11220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11219_3_lut (.I0(\mem_REG.mem_4_2 ), .I1(\mem_REG.mem_5_2 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13330));
    defparam i11219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_13381  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_29 ), .I2(\mem_REG.mem_3_29 ), .I3(rd_addr_r[1]), 
            .O(n15679));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_13381 .LUT_INIT = 16'he4aa;
    SB_LUT4 n15679_bdd_4_lut (.I0(n15679), .I1(\mem_REG.mem_1_29 ), .I2(\mem_REG.mem_0_29 ), 
            .I3(rd_addr_r[1]), .O(n15682));
    defparam n15679_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13406 (.I0(rd_addr_r[1]), .I1(n13777), 
            .I2(n13778), .I3(rd_addr_r[2]), .O(n15661));
    defparam rd_addr_r_1__bdd_4_lut_13406.LUT_INIT = 16'he4aa;
    SB_LUT4 n15661_bdd_4_lut (.I0(n15661), .I1(n13670), .I2(n13669), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[26]));
    defparam n15661_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11642_3_lut (.I0(\mem_REG.mem_0_25 ), .I1(\mem_REG.mem_1_25 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13753));
    defparam i11642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11643_3_lut (.I0(\mem_REG.mem_2_25 ), .I1(\mem_REG.mem_3_25 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13754));
    defparam i11643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11562_3_lut (.I0(\mem_REG.mem_6_25 ), .I1(\mem_REG.mem_7_25 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13673));
    defparam i11562_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11561_3_lut (.I0(\mem_REG.mem_4_25 ), .I1(\mem_REG.mem_5_25 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13672));
    defparam i11561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5371_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[31] ), 
            .I3(\mem_REG.mem_6_31 ), .O(n6845));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5371_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5370_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[30] ), 
            .I3(\mem_REG.mem_6_30 ), .O(n6844));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5370_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5369_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[29] ), 
            .I3(\mem_REG.mem_6_29 ), .O(n6843));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5369_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5368_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[28] ), 
            .I3(\mem_REG.mem_6_28 ), .O(n6842));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5368_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5367_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[27] ), 
            .I3(\mem_REG.mem_6_27 ), .O(n6841));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5367_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5366_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[26] ), 
            .I3(\mem_REG.mem_6_26 ), .O(n6840));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5366_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5365_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[25] ), 
            .I3(\mem_REG.mem_6_25 ), .O(n6839));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5365_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5364_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[24] ), 
            .I3(\mem_REG.mem_6_24 ), .O(n6838));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5364_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5363_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[23] ), 
            .I3(\mem_REG.mem_6_23 ), .O(n6837));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5363_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5362_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[22] ), 
            .I3(\mem_REG.mem_6_22 ), .O(n6836));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5362_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5361_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[21] ), 
            .I3(\mem_REG.mem_6_21 ), .O(n6835));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5361_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5360_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[20] ), 
            .I3(\mem_REG.mem_6_20 ), .O(n6834));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5360_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5359_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[19] ), 
            .I3(\mem_REG.mem_6_19 ), .O(n6833));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5359_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5358_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[18] ), 
            .I3(\mem_REG.mem_6_18 ), .O(n6832));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5358_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5357_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[17] ), 
            .I3(\mem_REG.mem_6_17 ), .O(n6831));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5357_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5356_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[16] ), 
            .I3(\mem_REG.mem_6_16 ), .O(n6830));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5356_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5355_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[15] ), 
            .I3(\mem_REG.mem_6_15 ), .O(n6829));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5355_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5354_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[14] ), 
            .I3(\mem_REG.mem_6_14 ), .O(n6828));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5354_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5353_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[13] ), 
            .I3(\mem_REG.mem_6_13 ), .O(n6827));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5353_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5352_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[12] ), 
            .I3(\mem_REG.mem_6_12 ), .O(n6826));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5352_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5351_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[11] ), 
            .I3(\mem_REG.mem_6_11 ), .O(n6825));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5351_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5350_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[10] ), 
            .I3(\mem_REG.mem_6_10 ), .O(n6824));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5350_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5349_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[9] ), 
            .I3(\mem_REG.mem_6_9 ), .O(n6823));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5349_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5348_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[8] ), 
            .I3(\mem_REG.mem_6_8 ), .O(n6822));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5348_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5347_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[7] ), 
            .I3(\mem_REG.mem_6_7 ), .O(n6821));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5347_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5346_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[6] ), 
            .I3(\mem_REG.mem_6_6 ), .O(n6820));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5346_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5345_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[5] ), 
            .I3(\mem_REG.mem_6_5 ), .O(n6819));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5345_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5344_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[4] ), 
            .I3(\mem_REG.mem_6_4 ), .O(n6818));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5344_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5343_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[3] ), 
            .I3(\mem_REG.mem_6_3 ), .O(n6817));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5343_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5342_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[2] ), 
            .I3(\mem_REG.mem_6_2 ), .O(n6816));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5342_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5341_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[1] ), 
            .I3(\mem_REG.mem_6_1 ), .O(n6815));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5341_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5340_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(DEBUG_5_c_0), 
            .I3(\mem_REG.mem_6_0 ), .O(n6814));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5340_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i803_804 (.Q(\mem_REG.mem_7_31 ), .C(SLM_CLK_c), .D(n6877));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i800_801 (.Q(\mem_REG.mem_7_30 ), .C(SLM_CLK_c), .D(n6876));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i797_798 (.Q(\mem_REG.mem_7_29 ), .C(SLM_CLK_c), .D(n6875));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i794_795 (.Q(\mem_REG.mem_7_28 ), .C(SLM_CLK_c), .D(n6874));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i791_792 (.Q(\mem_REG.mem_7_27 ), .C(SLM_CLK_c), .D(n6873));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i788_789 (.Q(\mem_REG.mem_7_26 ), .C(SLM_CLK_c), .D(n6872));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i785_786 (.Q(\mem_REG.mem_7_25 ), .C(SLM_CLK_c), .D(n6871));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i782_783 (.Q(\mem_REG.mem_7_24 ), .C(SLM_CLK_c), .D(n6870));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i779_780 (.Q(\mem_REG.mem_7_23 ), .C(SLM_CLK_c), .D(n6869));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i776_777 (.Q(\mem_REG.mem_7_22 ), .C(SLM_CLK_c), .D(n6868));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i773_774 (.Q(\mem_REG.mem_7_21 ), .C(SLM_CLK_c), .D(n6867));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i770_771 (.Q(\mem_REG.mem_7_20 ), .C(SLM_CLK_c), .D(n6866));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i767_768 (.Q(\mem_REG.mem_7_19 ), .C(SLM_CLK_c), .D(n6865));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i764_765 (.Q(\mem_REG.mem_7_18 ), .C(SLM_CLK_c), .D(n6864));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i761_762 (.Q(\mem_REG.mem_7_17 ), .C(SLM_CLK_c), .D(n6863));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i758_759 (.Q(\mem_REG.mem_7_16 ), .C(SLM_CLK_c), .D(n6862));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i755_756 (.Q(\mem_REG.mem_7_15 ), .C(SLM_CLK_c), .D(n6861));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i752_753 (.Q(\mem_REG.mem_7_14 ), .C(SLM_CLK_c), .D(n6860));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i749_750 (.Q(\mem_REG.mem_7_13 ), .C(SLM_CLK_c), .D(n6859));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i746_747 (.Q(\mem_REG.mem_7_12 ), .C(SLM_CLK_c), .D(n6858));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i743_744 (.Q(\mem_REG.mem_7_11 ), .C(SLM_CLK_c), .D(n6857));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i740_741 (.Q(\mem_REG.mem_7_10 ), .C(SLM_CLK_c), .D(n6856));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i737_738 (.Q(\mem_REG.mem_7_9 ), .C(SLM_CLK_c), .D(n6855));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i734_735 (.Q(\mem_REG.mem_7_8 ), .C(SLM_CLK_c), .D(n6854));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i731_732 (.Q(\mem_REG.mem_7_7 ), .C(SLM_CLK_c), .D(n6853));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i728_729 (.Q(\mem_REG.mem_7_6 ), .C(SLM_CLK_c), .D(n6852));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i725_726 (.Q(\mem_REG.mem_7_5 ), .C(SLM_CLK_c), .D(n6851));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i722_723 (.Q(\mem_REG.mem_7_4 ), .C(SLM_CLK_c), .D(n6850));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i719_720 (.Q(\mem_REG.mem_7_3 ), .C(SLM_CLK_c), .D(n6849));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i716_717 (.Q(\mem_REG.mem_7_2 ), .C(SLM_CLK_c), .D(n6848));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i713_714 (.Q(\mem_REG.mem_7_1 ), .C(SLM_CLK_c), .D(n6847));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i710_711 (.Q(\mem_REG.mem_7_0 ), .C(SLM_CLK_c), .D(n6846));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i707_708 (.Q(\mem_REG.mem_6_31 ), .C(SLM_CLK_c), .D(n6845));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i704_705 (.Q(\mem_REG.mem_6_30 ), .C(SLM_CLK_c), .D(n6844));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i701_702 (.Q(\mem_REG.mem_6_29 ), .C(SLM_CLK_c), .D(n6843));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i698_699 (.Q(\mem_REG.mem_6_28 ), .C(SLM_CLK_c), .D(n6842));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i695_696 (.Q(\mem_REG.mem_6_27 ), .C(SLM_CLK_c), .D(n6841));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i692_693 (.Q(\mem_REG.mem_6_26 ), .C(SLM_CLK_c), .D(n6840));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i689_690 (.Q(\mem_REG.mem_6_25 ), .C(SLM_CLK_c), .D(n6839));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i686_687 (.Q(\mem_REG.mem_6_24 ), .C(SLM_CLK_c), .D(n6838));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i683_684 (.Q(\mem_REG.mem_6_23 ), .C(SLM_CLK_c), .D(n6837));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i680_681 (.Q(\mem_REG.mem_6_22 ), .C(SLM_CLK_c), .D(n6836));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i677_678 (.Q(\mem_REG.mem_6_21 ), .C(SLM_CLK_c), .D(n6835));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i674_675 (.Q(\mem_REG.mem_6_20 ), .C(SLM_CLK_c), .D(n6834));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i671_672 (.Q(\mem_REG.mem_6_19 ), .C(SLM_CLK_c), .D(n6833));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i668_669 (.Q(\mem_REG.mem_6_18 ), .C(SLM_CLK_c), .D(n6832));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i665_666 (.Q(\mem_REG.mem_6_17 ), .C(SLM_CLK_c), .D(n6831));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i662_663 (.Q(\mem_REG.mem_6_16 ), .C(SLM_CLK_c), .D(n6830));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i659_660 (.Q(\mem_REG.mem_6_15 ), .C(SLM_CLK_c), .D(n6829));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i656_657 (.Q(\mem_REG.mem_6_14 ), .C(SLM_CLK_c), .D(n6828));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i653_654 (.Q(\mem_REG.mem_6_13 ), .C(SLM_CLK_c), .D(n6827));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i650_651 (.Q(\mem_REG.mem_6_12 ), .C(SLM_CLK_c), .D(n6826));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i647_648 (.Q(\mem_REG.mem_6_11 ), .C(SLM_CLK_c), .D(n6825));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i644_645 (.Q(\mem_REG.mem_6_10 ), .C(SLM_CLK_c), .D(n6824));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i641_642 (.Q(\mem_REG.mem_6_9 ), .C(SLM_CLK_c), .D(n6823));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i638_639 (.Q(\mem_REG.mem_6_8 ), .C(SLM_CLK_c), .D(n6822));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i635_636 (.Q(\mem_REG.mem_6_7 ), .C(SLM_CLK_c), .D(n6821));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i632_633 (.Q(\mem_REG.mem_6_6 ), .C(SLM_CLK_c), .D(n6820));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i629_630 (.Q(\mem_REG.mem_6_5 ), .C(SLM_CLK_c), .D(n6819));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i626_627 (.Q(\mem_REG.mem_6_4 ), .C(SLM_CLK_c), .D(n6818));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i623_624 (.Q(\mem_REG.mem_6_3 ), .C(SLM_CLK_c), .D(n6817));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i620_621 (.Q(\mem_REG.mem_6_2 ), .C(SLM_CLK_c), .D(n6816));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i617_618 (.Q(\mem_REG.mem_6_1 ), .C(SLM_CLK_c), .D(n6815));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i614_615 (.Q(\mem_REG.mem_6_0 ), .C(SLM_CLK_c), .D(n6814));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i611_612 (.Q(\mem_REG.mem_5_31 ), .C(SLM_CLK_c), .D(n6813));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i608_609 (.Q(\mem_REG.mem_5_30 ), .C(SLM_CLK_c), .D(n6812));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i605_606 (.Q(\mem_REG.mem_5_29 ), .C(SLM_CLK_c), .D(n6811));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i602_603 (.Q(\mem_REG.mem_5_28 ), .C(SLM_CLK_c), .D(n6810));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i599_600 (.Q(\mem_REG.mem_5_27 ), .C(SLM_CLK_c), .D(n6809));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i596_597 (.Q(\mem_REG.mem_5_26 ), .C(SLM_CLK_c), .D(n6808));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i593_594 (.Q(\mem_REG.mem_5_25 ), .C(SLM_CLK_c), .D(n6807));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i590_591 (.Q(\mem_REG.mem_5_24 ), .C(SLM_CLK_c), .D(n6806));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i587_588 (.Q(\mem_REG.mem_5_23 ), .C(SLM_CLK_c), .D(n6805));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i584_585 (.Q(\mem_REG.mem_5_22 ), .C(SLM_CLK_c), .D(n6804));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i581_582 (.Q(\mem_REG.mem_5_21 ), .C(SLM_CLK_c), .D(n6803));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i578_579 (.Q(\mem_REG.mem_5_20 ), .C(SLM_CLK_c), .D(n6802));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i575_576 (.Q(\mem_REG.mem_5_19 ), .C(SLM_CLK_c), .D(n6801));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i572_573 (.Q(\mem_REG.mem_5_18 ), .C(SLM_CLK_c), .D(n6800));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i569_570 (.Q(\mem_REG.mem_5_17 ), .C(SLM_CLK_c), .D(n6799));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i566_567 (.Q(\mem_REG.mem_5_16 ), .C(SLM_CLK_c), .D(n6798));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i563_564 (.Q(\mem_REG.mem_5_15 ), .C(SLM_CLK_c), .D(n6797));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i560_561 (.Q(\mem_REG.mem_5_14 ), .C(SLM_CLK_c), .D(n6796));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i557_558 (.Q(\mem_REG.mem_5_13 ), .C(SLM_CLK_c), .D(n6795));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i554_555 (.Q(\mem_REG.mem_5_12 ), .C(SLM_CLK_c), .D(n6794));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i551_552 (.Q(\mem_REG.mem_5_11 ), .C(SLM_CLK_c), .D(n6793));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i548_549 (.Q(\mem_REG.mem_5_10 ), .C(SLM_CLK_c), .D(n6792));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i545_546 (.Q(\mem_REG.mem_5_9 ), .C(SLM_CLK_c), .D(n6791));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i542_543 (.Q(\mem_REG.mem_5_8 ), .C(SLM_CLK_c), .D(n6790));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i539_540 (.Q(\mem_REG.mem_5_7 ), .C(SLM_CLK_c), .D(n6789));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i536_537 (.Q(\mem_REG.mem_5_6 ), .C(SLM_CLK_c), .D(n6788));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i533_534 (.Q(\mem_REG.mem_5_5 ), .C(SLM_CLK_c), .D(n6787));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i530_531 (.Q(\mem_REG.mem_5_4 ), .C(SLM_CLK_c), .D(n6786));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i527_528 (.Q(\mem_REG.mem_5_3 ), .C(SLM_CLK_c), .D(n6785));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i524_525 (.Q(\mem_REG.mem_5_2 ), .C(SLM_CLK_c), .D(n6784));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i521_522 (.Q(\mem_REG.mem_5_1 ), .C(SLM_CLK_c), .D(n6783));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i518_519 (.Q(\mem_REG.mem_5_0 ), .C(SLM_CLK_c), .D(n6782));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i515_516 (.Q(\mem_REG.mem_4_31 ), .C(SLM_CLK_c), .D(n6781));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i512_513 (.Q(\mem_REG.mem_4_30 ), .C(SLM_CLK_c), .D(n6780));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i509_510 (.Q(\mem_REG.mem_4_29 ), .C(SLM_CLK_c), .D(n6779));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i506_507 (.Q(\mem_REG.mem_4_28 ), .C(SLM_CLK_c), .D(n6778));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i503_504 (.Q(\mem_REG.mem_4_27 ), .C(SLM_CLK_c), .D(n6777));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i500_501 (.Q(\mem_REG.mem_4_26 ), .C(SLM_CLK_c), .D(n6776));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i497_498 (.Q(\mem_REG.mem_4_25 ), .C(SLM_CLK_c), .D(n6775));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i494_495 (.Q(\mem_REG.mem_4_24 ), .C(SLM_CLK_c), .D(n6774));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i491_492 (.Q(\mem_REG.mem_4_23 ), .C(SLM_CLK_c), .D(n6773));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i488_489 (.Q(\mem_REG.mem_4_22 ), .C(SLM_CLK_c), .D(n6772));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i485_486 (.Q(\mem_REG.mem_4_21 ), .C(SLM_CLK_c), .D(n6771));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i482_483 (.Q(\mem_REG.mem_4_20 ), .C(SLM_CLK_c), .D(n6770));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i479_480 (.Q(\mem_REG.mem_4_19 ), .C(SLM_CLK_c), .D(n6769));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i476_477 (.Q(\mem_REG.mem_4_18 ), .C(SLM_CLK_c), .D(n6768));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i473_474 (.Q(\mem_REG.mem_4_17 ), .C(SLM_CLK_c), .D(n6767));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i470_471 (.Q(\mem_REG.mem_4_16 ), .C(SLM_CLK_c), .D(n6766));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i467_468 (.Q(\mem_REG.mem_4_15 ), .C(SLM_CLK_c), .D(n6765));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i464_465 (.Q(\mem_REG.mem_4_14 ), .C(SLM_CLK_c), .D(n6764));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i461_462 (.Q(\mem_REG.mem_4_13 ), .C(SLM_CLK_c), .D(n6763));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i458_459 (.Q(\mem_REG.mem_4_12 ), .C(SLM_CLK_c), .D(n6762));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i455_456 (.Q(\mem_REG.mem_4_11 ), .C(SLM_CLK_c), .D(n6761));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i452_453 (.Q(\mem_REG.mem_4_10 ), .C(SLM_CLK_c), .D(n6760));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i449_450 (.Q(\mem_REG.mem_4_9 ), .C(SLM_CLK_c), .D(n6759));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i446_447 (.Q(\mem_REG.mem_4_8 ), .C(SLM_CLK_c), .D(n6758));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i443_444 (.Q(\mem_REG.mem_4_7 ), .C(SLM_CLK_c), .D(n6757));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i440_441 (.Q(\mem_REG.mem_4_6 ), .C(SLM_CLK_c), .D(n6756));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i437_438 (.Q(\mem_REG.mem_4_5 ), .C(SLM_CLK_c), .D(n6755));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i434_435 (.Q(\mem_REG.mem_4_4 ), .C(SLM_CLK_c), .D(n6754));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i431_432 (.Q(\mem_REG.mem_4_3 ), .C(SLM_CLK_c), .D(n6753));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i428_429 (.Q(\mem_REG.mem_4_2 ), .C(SLM_CLK_c), .D(n6752));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i425_426 (.Q(\mem_REG.mem_4_1 ), .C(SLM_CLK_c), .D(n6751));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i422_423 (.Q(\mem_REG.mem_4_0 ), .C(SLM_CLK_c), .D(n6750));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i419_420 (.Q(\mem_REG.mem_3_31 ), .C(SLM_CLK_c), .D(n6749));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i416_417 (.Q(\mem_REG.mem_3_30 ), .C(SLM_CLK_c), .D(n6748));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i413_414 (.Q(\mem_REG.mem_3_29 ), .C(SLM_CLK_c), .D(n6747));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i410_411 (.Q(\mem_REG.mem_3_28 ), .C(SLM_CLK_c), .D(n6746));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i407_408 (.Q(\mem_REG.mem_3_27 ), .C(SLM_CLK_c), .D(n6745));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i404_405 (.Q(\mem_REG.mem_3_26 ), .C(SLM_CLK_c), .D(n6744));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i401_402 (.Q(\mem_REG.mem_3_25 ), .C(SLM_CLK_c), .D(n6743));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i398_399 (.Q(\mem_REG.mem_3_24 ), .C(SLM_CLK_c), .D(n6742));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i395_396 (.Q(\mem_REG.mem_3_23 ), .C(SLM_CLK_c), .D(n6741));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i392_393 (.Q(\mem_REG.mem_3_22 ), .C(SLM_CLK_c), .D(n6740));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i389_390 (.Q(\mem_REG.mem_3_21 ), .C(SLM_CLK_c), .D(n6739));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i386_387 (.Q(\mem_REG.mem_3_20 ), .C(SLM_CLK_c), .D(n6738));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i383_384 (.Q(\mem_REG.mem_3_19 ), .C(SLM_CLK_c), .D(n6737));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i380_381 (.Q(\mem_REG.mem_3_18 ), .C(SLM_CLK_c), .D(n6736));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i377_378 (.Q(\mem_REG.mem_3_17 ), .C(SLM_CLK_c), .D(n6735));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i374_375 (.Q(\mem_REG.mem_3_16 ), .C(SLM_CLK_c), .D(n6734));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i371_372 (.Q(\mem_REG.mem_3_15 ), .C(SLM_CLK_c), .D(n6733));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i368_369 (.Q(\mem_REG.mem_3_14 ), .C(SLM_CLK_c), .D(n6732));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i365_366 (.Q(\mem_REG.mem_3_13 ), .C(SLM_CLK_c), .D(n6731));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i362_363 (.Q(\mem_REG.mem_3_12 ), .C(SLM_CLK_c), .D(n6730));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i359_360 (.Q(\mem_REG.mem_3_11 ), .C(SLM_CLK_c), .D(n6729));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i356_357 (.Q(\mem_REG.mem_3_10 ), .C(SLM_CLK_c), .D(n6728));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i353_354 (.Q(\mem_REG.mem_3_9 ), .C(SLM_CLK_c), .D(n6727));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i350_351 (.Q(\mem_REG.mem_3_8 ), .C(SLM_CLK_c), .D(n6726));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i347_348 (.Q(\mem_REG.mem_3_7 ), .C(SLM_CLK_c), .D(n6725));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i344_345 (.Q(\mem_REG.mem_3_6 ), .C(SLM_CLK_c), .D(n6724));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i341_342 (.Q(\mem_REG.mem_3_5 ), .C(SLM_CLK_c), .D(n6723));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i338_339 (.Q(\mem_REG.mem_3_4 ), .C(SLM_CLK_c), .D(n6722));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i335_336 (.Q(\mem_REG.mem_3_3 ), .C(SLM_CLK_c), .D(n6721));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i332_333 (.Q(\mem_REG.mem_3_2 ), .C(SLM_CLK_c), .D(n6720));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i329_330 (.Q(\mem_REG.mem_3_1 ), .C(SLM_CLK_c), .D(n6719));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i326_327 (.Q(\mem_REG.mem_3_0 ), .C(SLM_CLK_c), .D(n6718));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i323_324 (.Q(\mem_REG.mem_2_31 ), .C(SLM_CLK_c), .D(n6717));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i320_321 (.Q(\mem_REG.mem_2_30 ), .C(SLM_CLK_c), .D(n6716));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i317_318 (.Q(\mem_REG.mem_2_29 ), .C(SLM_CLK_c), .D(n6715));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i314_315 (.Q(\mem_REG.mem_2_28 ), .C(SLM_CLK_c), .D(n6714));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i311_312 (.Q(\mem_REG.mem_2_27 ), .C(SLM_CLK_c), .D(n6713));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i308_309 (.Q(\mem_REG.mem_2_26 ), .C(SLM_CLK_c), .D(n6712));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i305_306 (.Q(\mem_REG.mem_2_25 ), .C(SLM_CLK_c), .D(n6711));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i302_303 (.Q(\mem_REG.mem_2_24 ), .C(SLM_CLK_c), .D(n6710));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i299_300 (.Q(\mem_REG.mem_2_23 ), .C(SLM_CLK_c), .D(n6709));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i296_297 (.Q(\mem_REG.mem_2_22 ), .C(SLM_CLK_c), .D(n6708));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i293_294 (.Q(\mem_REG.mem_2_21 ), .C(SLM_CLK_c), .D(n6707));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i290_291 (.Q(\mem_REG.mem_2_20 ), .C(SLM_CLK_c), .D(n6706));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i287_288 (.Q(\mem_REG.mem_2_19 ), .C(SLM_CLK_c), .D(n6705));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i284_285 (.Q(\mem_REG.mem_2_18 ), .C(SLM_CLK_c), .D(n6704));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i281_282 (.Q(\mem_REG.mem_2_17 ), .C(SLM_CLK_c), .D(n6703));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i278_279 (.Q(\mem_REG.mem_2_16 ), .C(SLM_CLK_c), .D(n6702));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i275_276 (.Q(\mem_REG.mem_2_15 ), .C(SLM_CLK_c), .D(n6701));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i272_273 (.Q(\mem_REG.mem_2_14 ), .C(SLM_CLK_c), .D(n6700));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i269_270 (.Q(\mem_REG.mem_2_13 ), .C(SLM_CLK_c), .D(n6699));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i266_267 (.Q(\mem_REG.mem_2_12 ), .C(SLM_CLK_c), .D(n6698));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i263_264 (.Q(\mem_REG.mem_2_11 ), .C(SLM_CLK_c), .D(n6697));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i260_261 (.Q(\mem_REG.mem_2_10 ), .C(SLM_CLK_c), .D(n6696));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i257_258 (.Q(\mem_REG.mem_2_9 ), .C(SLM_CLK_c), .D(n6695));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i254_255 (.Q(\mem_REG.mem_2_8 ), .C(SLM_CLK_c), .D(n6694));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i251_252 (.Q(\mem_REG.mem_2_7 ), .C(SLM_CLK_c), .D(n6693));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i248_249 (.Q(\mem_REG.mem_2_6 ), .C(SLM_CLK_c), .D(n6692));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i245_246 (.Q(\mem_REG.mem_2_5 ), .C(SLM_CLK_c), .D(n6691));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i242_243 (.Q(\mem_REG.mem_2_4 ), .C(SLM_CLK_c), .D(n6690));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i239_240 (.Q(\mem_REG.mem_2_3 ), .C(SLM_CLK_c), .D(n6689));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i236_237 (.Q(\mem_REG.mem_2_2 ), .C(SLM_CLK_c), .D(n6688));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i233_234 (.Q(\mem_REG.mem_2_1 ), .C(SLM_CLK_c), .D(n6687));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i230_231 (.Q(\mem_REG.mem_2_0 ), .C(SLM_CLK_c), .D(n6686));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i227_228 (.Q(\mem_REG.mem_1_31 ), .C(SLM_CLK_c), .D(n6685));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i224_225 (.Q(\mem_REG.mem_1_30 ), .C(SLM_CLK_c), .D(n6684));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i221_222 (.Q(\mem_REG.mem_1_29 ), .C(SLM_CLK_c), .D(n6683));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i218_219 (.Q(\mem_REG.mem_1_28 ), .C(SLM_CLK_c), .D(n6682));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i215_216 (.Q(\mem_REG.mem_1_27 ), .C(SLM_CLK_c), .D(n6681));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i212_213 (.Q(\mem_REG.mem_1_26 ), .C(SLM_CLK_c), .D(n6680));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i209_210 (.Q(\mem_REG.mem_1_25 ), .C(SLM_CLK_c), .D(n6679));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i206_207 (.Q(\mem_REG.mem_1_24 ), .C(SLM_CLK_c), .D(n6678));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i203_204 (.Q(\mem_REG.mem_1_23 ), .C(SLM_CLK_c), .D(n6677));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i200_201 (.Q(\mem_REG.mem_1_22 ), .C(SLM_CLK_c), .D(n6676));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i197_198 (.Q(\mem_REG.mem_1_21 ), .C(SLM_CLK_c), .D(n6675));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i194_195 (.Q(\mem_REG.mem_1_20 ), .C(SLM_CLK_c), .D(n6674));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i191_192 (.Q(\mem_REG.mem_1_19 ), .C(SLM_CLK_c), .D(n6673));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i188_189 (.Q(\mem_REG.mem_1_18 ), .C(SLM_CLK_c), .D(n6672));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i185_186 (.Q(\mem_REG.mem_1_17 ), .C(SLM_CLK_c), .D(n6671));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i182_183 (.Q(\mem_REG.mem_1_16 ), .C(SLM_CLK_c), .D(n6670));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i179_180 (.Q(\mem_REG.mem_1_15 ), .C(SLM_CLK_c), .D(n6669));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i176_177 (.Q(\mem_REG.mem_1_14 ), .C(SLM_CLK_c), .D(n6668));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i173_174 (.Q(\mem_REG.mem_1_13 ), .C(SLM_CLK_c), .D(n6667));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i170_171 (.Q(\mem_REG.mem_1_12 ), .C(SLM_CLK_c), .D(n6666));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i167_168 (.Q(\mem_REG.mem_1_11 ), .C(SLM_CLK_c), .D(n6665));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i164_165 (.Q(\mem_REG.mem_1_10 ), .C(SLM_CLK_c), .D(n6664));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i161_162 (.Q(\mem_REG.mem_1_9 ), .C(SLM_CLK_c), .D(n6663));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i158_159 (.Q(\mem_REG.mem_1_8 ), .C(SLM_CLK_c), .D(n6662));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i155_156 (.Q(\mem_REG.mem_1_7 ), .C(SLM_CLK_c), .D(n6661));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i152_153 (.Q(\mem_REG.mem_1_6 ), .C(SLM_CLK_c), .D(n6660));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i149_150 (.Q(\mem_REG.mem_1_5 ), .C(SLM_CLK_c), .D(n6659));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i146_147 (.Q(\mem_REG.mem_1_4 ), .C(SLM_CLK_c), .D(n6658));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i143_144 (.Q(\mem_REG.mem_1_3 ), .C(SLM_CLK_c), .D(n6657));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i140_141 (.Q(\mem_REG.mem_1_2 ), .C(SLM_CLK_c), .D(n6656));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i137_138 (.Q(\mem_REG.mem_1_1 ), .C(SLM_CLK_c), .D(n6655));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i134_135 (.Q(\mem_REG.mem_1_0 ), .C(SLM_CLK_c), .D(n6654));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i131_132 (.Q(\mem_REG.mem_0_31 ), .C(SLM_CLK_c), .D(n6653));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i128_129 (.Q(\mem_REG.mem_0_30 ), .C(SLM_CLK_c), .D(n6652));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i125_126 (.Q(\mem_REG.mem_0_29 ), .C(SLM_CLK_c), .D(n6651));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i122_123 (.Q(\mem_REG.mem_0_28 ), .C(SLM_CLK_c), .D(n6650));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i119_120 (.Q(\mem_REG.mem_0_27 ), .C(SLM_CLK_c), .D(n6649));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i116_117 (.Q(\mem_REG.mem_0_26 ), .C(SLM_CLK_c), .D(n6648));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i113_114 (.Q(\mem_REG.mem_0_25 ), .C(SLM_CLK_c), .D(n6647));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i110_111 (.Q(\mem_REG.mem_0_24 ), .C(SLM_CLK_c), .D(n6646));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i107_108 (.Q(\mem_REG.mem_0_23 ), .C(SLM_CLK_c), .D(n6645));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i104_105 (.Q(\mem_REG.mem_0_22 ), .C(SLM_CLK_c), .D(n6644));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i101_102 (.Q(\mem_REG.mem_0_21 ), .C(SLM_CLK_c), .D(n6643));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i98_99 (.Q(\mem_REG.mem_0_20 ), .C(SLM_CLK_c), .D(n6642));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i95_96 (.Q(\mem_REG.mem_0_19 ), .C(SLM_CLK_c), .D(n6641));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i92_93 (.Q(\mem_REG.mem_0_18 ), .C(SLM_CLK_c), .D(n6640));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i89_90 (.Q(\mem_REG.mem_0_17 ), .C(SLM_CLK_c), .D(n6639));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i86_87 (.Q(\mem_REG.mem_0_16 ), .C(SLM_CLK_c), .D(n6638));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i83_84 (.Q(\mem_REG.mem_0_15 ), .C(SLM_CLK_c), .D(n6637));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i80_81 (.Q(\mem_REG.mem_0_14 ), .C(SLM_CLK_c), .D(n6636));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i77_78 (.Q(\mem_REG.mem_0_13 ), .C(SLM_CLK_c), .D(n6635));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i74_75 (.Q(\mem_REG.mem_0_12 ), .C(SLM_CLK_c), .D(n6634));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i71_72 (.Q(\mem_REG.mem_0_11 ), .C(SLM_CLK_c), .D(n6633));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i68_69 (.Q(\mem_REG.mem_0_10 ), .C(SLM_CLK_c), .D(n6632));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i65_66 (.Q(\mem_REG.mem_0_9 ), .C(SLM_CLK_c), .D(n6631));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i62_63 (.Q(\mem_REG.mem_0_8 ), .C(SLM_CLK_c), .D(n6630));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i59_60 (.Q(\mem_REG.mem_0_7 ), .C(SLM_CLK_c), .D(n6629));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i56_57 (.Q(\mem_REG.mem_0_6 ), .C(SLM_CLK_c), .D(n6628));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i53_54 (.Q(\mem_REG.mem_0_5 ), .C(SLM_CLK_c), .D(n6627));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i50_51 (.Q(\mem_REG.mem_0_4 ), .C(SLM_CLK_c), .D(n6626));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i47_48 (.Q(\mem_REG.mem_0_3 ), .C(SLM_CLK_c), .D(n6625));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i44_45 (.Q(\mem_REG.mem_0_2 ), .C(SLM_CLK_c), .D(n6624));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i41_42 (.Q(\mem_REG.mem_0_1 ), .C(SLM_CLK_c), .D(n6623));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i38_39 (.Q(\mem_REG.mem_0_0 ), .C(SLM_CLK_c), .D(n6622));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_LUT4 i11558_3_lut (.I0(\mem_REG.mem_0_26 ), .I1(\mem_REG.mem_1_26 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13669));
    defparam i11558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11559_3_lut (.I0(\mem_REG.mem_2_26 ), .I1(\mem_REG.mem_3_26 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13670));
    defparam i11559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13351 (.I0(rd_addr_r[1]), .I1(n13672), 
            .I2(n13673), .I3(rd_addr_r[2]), .O(n15619));
    defparam rd_addr_r_1__bdd_4_lut_13351.LUT_INIT = 16'he4aa;
    SB_LUT4 n15619_bdd_4_lut (.I0(n15619), .I1(n13754), .I2(n13753), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[25]));
    defparam n15619_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5339_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[31] ), 
            .I3(\mem_REG.mem_5_31 ), .O(n6813));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5339_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5338_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[30] ), 
            .I3(\mem_REG.mem_5_30 ), .O(n6812));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5338_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5337_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[29] ), 
            .I3(\mem_REG.mem_5_29 ), .O(n6811));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5337_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5336_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[28] ), 
            .I3(\mem_REG.mem_5_28 ), .O(n6810));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5336_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11667_3_lut (.I0(\mem_REG.mem_6_26 ), .I1(\mem_REG.mem_7_26 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13778));
    defparam i11667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5335_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[27] ), 
            .I3(\mem_REG.mem_5_27 ), .O(n6809));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5335_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11666_3_lut (.I0(\mem_REG.mem_4_26 ), .I1(\mem_REG.mem_5_26 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13777));
    defparam i11666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5334_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[26] ), 
            .I3(\mem_REG.mem_5_26 ), .O(n6808));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5334_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5333_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[25] ), 
            .I3(\mem_REG.mem_5_25 ), .O(n6807));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5333_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5332_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[24] ), 
            .I3(\mem_REG.mem_5_24 ), .O(n6806));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5332_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5331_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[23] ), 
            .I3(\mem_REG.mem_5_23 ), .O(n6805));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5331_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5330_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[22] ), 
            .I3(\mem_REG.mem_5_22 ), .O(n6804));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5330_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5329_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[21] ), 
            .I3(\mem_REG.mem_5_21 ), .O(n6803));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5329_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5328_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[20] ), 
            .I3(\mem_REG.mem_5_20 ), .O(n6802));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5328_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5327_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[19] ), 
            .I3(\mem_REG.mem_5_19 ), .O(n6801));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5327_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5326_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[18] ), 
            .I3(\mem_REG.mem_5_18 ), .O(n6800));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5326_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5325_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[17] ), 
            .I3(\mem_REG.mem_5_17 ), .O(n6799));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5325_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5324_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[16] ), 
            .I3(\mem_REG.mem_5_16 ), .O(n6798));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5324_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5323_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[15] ), 
            .I3(\mem_REG.mem_5_15 ), .O(n6797));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5323_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5322_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[14] ), 
            .I3(\mem_REG.mem_5_14 ), .O(n6796));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5322_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5321_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[13] ), 
            .I3(\mem_REG.mem_5_13 ), .O(n6795));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5321_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5320_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[12] ), 
            .I3(\mem_REG.mem_5_12 ), .O(n6794));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5320_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5319_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[11] ), 
            .I3(\mem_REG.mem_5_11 ), .O(n6793));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5319_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5318_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[10] ), 
            .I3(\mem_REG.mem_5_10 ), .O(n6792));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5318_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5317_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[9] ), 
            .I3(\mem_REG.mem_5_9 ), .O(n6791));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5317_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5316_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[8] ), 
            .I3(\mem_REG.mem_5_8 ), .O(n6790));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5316_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5315_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[7] ), 
            .I3(\mem_REG.mem_5_7 ), .O(n6789));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5315_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_12443  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_4 ), .I2(\mem_REG.mem_7_4 ), .I3(rd_addr_r[1]), 
            .O(n14509));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_12443 .LUT_INIT = 16'he4aa;
    SB_LUT4 i5314_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[6] ), 
            .I3(\mem_REG.mem_5_6 ), .O(n6788));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5314_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5313_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[5] ), 
            .I3(\mem_REG.mem_5_5 ), .O(n6787));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5313_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_12498  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_13 ), .I2(\mem_REG.mem_7_13 ), .I3(rd_addr_r[1]), 
            .O(n14605));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_12498 .LUT_INIT = 16'he4aa;
    SB_LUT4 i5312_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[4] ), 
            .I3(\mem_REG.mem_5_4 ), .O(n6786));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5312_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5311_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[3] ), 
            .I3(\mem_REG.mem_5_3 ), .O(n6785));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5311_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5310_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[2] ), 
            .I3(\mem_REG.mem_5_2 ), .O(n6784));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5310_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5309_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[1] ), 
            .I3(\mem_REG.mem_5_1 ), .O(n6783));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5309_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5308_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(DEBUG_5_c_0), 
            .I3(\mem_REG.mem_5_0 ), .O(n6782));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5308_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5307_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[31] ), 
            .I3(\mem_REG.mem_4_31 ), .O(n6781));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5307_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5306_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[30] ), 
            .I3(\mem_REG.mem_4_30 ), .O(n6780));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5306_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5305_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[29] ), 
            .I3(\mem_REG.mem_4_29 ), .O(n6779));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5305_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5304_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[28] ), 
            .I3(\mem_REG.mem_4_28 ), .O(n6778));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5304_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5303_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[27] ), 
            .I3(\mem_REG.mem_4_27 ), .O(n6777));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5303_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14605_bdd_4_lut (.I0(n14605), .I1(\mem_REG.mem_5_13 ), .I2(\mem_REG.mem_4_13 ), 
            .I3(rd_addr_r[1]), .O(n14608));
    defparam n14605_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5302_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[26] ), 
            .I3(\mem_REG.mem_4_26 ), .O(n6776));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5302_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12787 (.I0(rd_addr_r[1]), .I1(n13330), 
            .I2(n13331), .I3(rd_addr_r[2]), .O(n14905));
    defparam rd_addr_r_1__bdd_4_lut_12787.LUT_INIT = 16'he4aa;
    SB_LUT4 n14905_bdd_4_lut (.I0(n14905), .I1(n13328), .I2(n13327), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[2]));
    defparam n14905_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5301_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[25] ), 
            .I3(\mem_REG.mem_4_25 ), .O(n6775));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5301_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5300_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[24] ), 
            .I3(\mem_REG.mem_4_24 ), .O(n6774));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5300_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5299_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[23] ), 
            .I3(\mem_REG.mem_4_23 ), .O(n6773));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5299_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5298_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[22] ), 
            .I3(\mem_REG.mem_4_22 ), .O(n6772));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5298_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5297_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[21] ), 
            .I3(\mem_REG.mem_4_21 ), .O(n6771));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5297_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13316 (.I0(rd_addr_r[1]), .I1(n13804), 
            .I2(n13805), .I3(rd_addr_r[2]), .O(n15589));
    defparam rd_addr_r_1__bdd_4_lut_13316.LUT_INIT = 16'he4aa;
    SB_LUT4 i5296_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[20] ), 
            .I3(\mem_REG.mem_4_20 ), .O(n6770));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5296_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5295_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[19] ), 
            .I3(\mem_REG.mem_4_19 ), .O(n6769));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5295_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5294_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[18] ), 
            .I3(\mem_REG.mem_4_18 ), .O(n6768));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5294_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5293_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[17] ), 
            .I3(\mem_REG.mem_4_17 ), .O(n6767));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5293_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15589_bdd_4_lut (.I0(n15589), .I1(n13745), .I2(n13744), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[9]));
    defparam n15589_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5292_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[16] ), 
            .I3(\mem_REG.mem_4_16 ), .O(n6766));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5292_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5291_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[15] ), 
            .I3(\mem_REG.mem_4_15 ), .O(n6765));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5291_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5290_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[14] ), 
            .I3(\mem_REG.mem_4_14 ), .O(n6764));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5290_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5289_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[13] ), 
            .I3(\mem_REG.mem_4_13 ), .O(n6763));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5289_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5288_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[12] ), 
            .I3(\mem_REG.mem_4_12 ), .O(n6762));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5288_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14509_bdd_4_lut (.I0(n14509), .I1(\mem_REG.mem_5_4 ), .I2(\mem_REG.mem_4_4 ), 
            .I3(rd_addr_r[1]), .O(n14512));
    defparam n14509_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5287_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[11] ), 
            .I3(\mem_REG.mem_4_11 ), .O(n6761));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5287_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5286_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[10] ), 
            .I3(\mem_REG.mem_4_10 ), .O(n6760));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5286_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5285_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[9] ), 
            .I3(\mem_REG.mem_4_9 ), .O(n6759));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5285_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5284_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[8] ), 
            .I3(\mem_REG.mem_4_8 ), .O(n6758));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5284_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13291 (.I0(rd_addr_r[1]), .I1(n13726), 
            .I2(n13727), .I3(rd_addr_r[2]), .O(n15577));
    defparam rd_addr_r_1__bdd_4_lut_13291.LUT_INIT = 16'he4aa;
    SB_LUT4 i5283_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[7] ), 
            .I3(\mem_REG.mem_4_7 ), .O(n6757));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5283_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n15577_bdd_4_lut (.I0(n15577), .I1(n13721), .I2(n13720), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[24]));
    defparam n15577_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5282_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[6] ), 
            .I3(\mem_REG.mem_4_6 ), .O(n6756));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5282_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5281_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[5] ), 
            .I3(\mem_REG.mem_4_5 ), .O(n6755));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5281_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5280_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[4] ), 
            .I3(\mem_REG.mem_4_4 ), .O(n6754));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5280_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5279_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[3] ), 
            .I3(\mem_REG.mem_4_3 ), .O(n6753));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5279_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5278_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[2] ), 
            .I3(\mem_REG.mem_4_2 ), .O(n6752));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5278_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5277_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[1] ), 
            .I3(\mem_REG.mem_4_1 ), .O(n6751));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5277_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5276_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(DEBUG_5_c_0), 
            .I3(\mem_REG.mem_4_0 ), .O(n6750));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5276_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13281 (.I0(rd_addr_r[1]), .I1(n13708), 
            .I2(n13709), .I3(rd_addr_r[2]), .O(n15559));
    defparam rd_addr_r_1__bdd_4_lut_13281.LUT_INIT = 16'he4aa;
    SB_LUT4 n15559_bdd_4_lut (.I0(n15559), .I1(n13679), .I2(n13678), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[8]));
    defparam n15559_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11039_3_lut (.I0(\mem_REG.mem_0_18 ), .I1(\mem_REG.mem_1_18 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13150));
    defparam i11039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11040_3_lut (.I0(\mem_REG.mem_2_18 ), .I1(\mem_REG.mem_3_18 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13151));
    defparam i11040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11622_3_lut (.I0(\mem_REG.mem_6_18 ), .I1(\mem_REG.mem_7_18 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13733));
    defparam i11622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11621_3_lut (.I0(\mem_REG.mem_4_18 ), .I1(\mem_REG.mem_5_18 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13732));
    defparam i11621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11318_3_lut (.I0(\mem_REG.mem_0_19 ), .I1(\mem_REG.mem_1_19 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13429));
    defparam i11318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11319_3_lut (.I0(\mem_REG.mem_2_19 ), .I1(\mem_REG.mem_3_19 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13430));
    defparam i11319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5275_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[31] ), 
            .I3(\mem_REG.mem_3_31 ), .O(n6749));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5275_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5274_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[30] ), 
            .I3(\mem_REG.mem_3_30 ), .O(n6748));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5274_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5273_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[29] ), 
            .I3(\mem_REG.mem_3_29 ), .O(n6747));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5273_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5272_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[28] ), 
            .I3(\mem_REG.mem_3_28 ), .O(n6746));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5272_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5271_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[27] ), 
            .I3(\mem_REG.mem_3_27 ), .O(n6745));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5271_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11613_3_lut (.I0(\mem_REG.mem_6_19 ), .I1(\mem_REG.mem_7_19 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13724));
    defparam i11613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5270_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[26] ), 
            .I3(\mem_REG.mem_3_26 ), .O(n6744));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5270_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11612_3_lut (.I0(\mem_REG.mem_4_19 ), .I1(\mem_REG.mem_5_19 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13723));
    defparam i11612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5269_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[25] ), 
            .I3(\mem_REG.mem_3_25 ), .O(n6743));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5269_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5268_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[24] ), 
            .I3(\mem_REG.mem_3_24 ), .O(n6742));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5268_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5267_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[23] ), 
            .I3(\mem_REG.mem_3_23 ), .O(n6741));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5267_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5266_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[22] ), 
            .I3(\mem_REG.mem_3_22 ), .O(n6740));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5266_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5265_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[21] ), 
            .I3(\mem_REG.mem_3_21 ), .O(n6739));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5265_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5264_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[20] ), 
            .I3(\mem_REG.mem_3_20 ), .O(n6738));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5264_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5263_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[19] ), 
            .I3(\mem_REG.mem_3_19 ), .O(n6737));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5263_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5262_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[18] ), 
            .I3(\mem_REG.mem_3_18 ), .O(n6736));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5262_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5261_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[17] ), 
            .I3(\mem_REG.mem_3_17 ), .O(n6735));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5261_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5260_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[16] ), 
            .I3(\mem_REG.mem_3_16 ), .O(n6734));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5260_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5259_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[15] ), 
            .I3(\mem_REG.mem_3_15 ), .O(n6733));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5259_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5258_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[14] ), 
            .I3(\mem_REG.mem_3_14 ), .O(n6732));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5258_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2221_3_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1cmp_r[2]), .I2(n3679), 
            .I3(GND_net), .O(n3402));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i2221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5257_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[13] ), 
            .I3(\mem_REG.mem_3_13 ), .O(n6731));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5257_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1751_3_lut (.I0(n2775[1]), .I1(n3400), .I2(n2), .I3(GND_net), 
            .O(n4));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i1751_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13266 (.I0(rd_addr_r[1]), .I1(n13687), 
            .I2(n13688), .I3(rd_addr_r[2]), .O(n15499));
    defparam rd_addr_r_1__bdd_4_lut_13266.LUT_INIT = 16'he4aa;
    SB_LUT4 i5256_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[12] ), 
            .I3(\mem_REG.mem_3_12 ), .O(n6730));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5256_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5255_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[11] ), 
            .I3(\mem_REG.mem_3_11 ), .O(n6729));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5255_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2219_3_lut (.I0(rd_addr_r[1]), .I1(rd_addr_p1cmp_r[1]), .I2(n3679), 
            .I3(GND_net), .O(n3400));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i2219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2044_3_lut (.I0(\MISC.rd_flag_addr_r [0]), .I1(\MISC.rd_flag_addr_p1_r [0]), 
            .I2(n3679), .I3(GND_net), .O(n3398));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i2044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1743_4_lut (.I0(\MISC.wr_flag_addr_r [0]), .I1(n3398), .I2(\MISC.wr_flag_addr_p1_r [0]), 
            .I3(n2057), .O(n2));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i1743_4_lut.LUT_INIT = 16'hf3bb;
    SB_LUT4 n15499_bdd_4_lut (.I0(n15499), .I1(n13676), .I2(n13675), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[22]));
    defparam n15499_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5254_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[10] ), 
            .I3(\mem_REG.mem_3_10 ), .O(n6728));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5254_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut (.I0(n2), .I1(n3400), .I2(n2775[1]), .I3(GND_net), 
            .O(n12302));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13216 (.I0(rd_addr_r[1]), .I1(n13714), 
            .I2(n13715), .I3(rd_addr_r[2]), .O(n15475));
    defparam rd_addr_r_1__bdd_4_lut_13216.LUT_INIT = 16'he4aa;
    SB_LUT4 i5253_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[9] ), 
            .I3(\mem_REG.mem_3_9 ), .O(n6727));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5253_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5252_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[8] ), 
            .I3(\mem_REG.mem_3_8 ), .O(n6726));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5252_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut (.I0(rd_addr_r[3]), .I1(n2775[3]), .I2(rd_addr_p1cmp_r[3]), 
            .I3(n3679), .O(n4_adj_1365));
    defparam i1_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_12473  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_4 ), .I2(\mem_REG.mem_3_4 ), .I3(rd_addr_r[1]), 
            .O(n14587));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_12473 .LUT_INIT = 16'he4aa;
    SB_LUT4 i5251_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[7] ), 
            .I3(\mem_REG.mem_3_7 ), .O(n6725));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5251_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_61 (.I0(n4), .I1(n3402), .I2(n2775[2]), .I3(GND_net), 
            .O(n12301));
    defparam i2_3_lut_adj_61.LUT_INIT = 16'h9696;
    SB_LUT4 i1758_3_lut (.I0(n2775[2]), .I1(n3402), .I2(n4), .I3(GND_net), 
            .O(n6_adj_1366));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i1758_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i2_4_lut (.I0(n6_adj_1366), .I1(n12301), .I2(n4_adj_1365), 
            .I3(n12302), .O(\MISC.AEmpty.almost_empty_nxt_w ));
    defparam i2_4_lut.LUT_INIT = 16'h4800;
    SB_LUT4 i10861_4_lut (.I0(rd_addr_p1cmp_r[1]), .I1(\MISC.rd_flag_addr_p1_r [0]), 
            .I2(wr_addr_r[1]), .I3(\MISC.wr_flag_addr_r [0]), .O(n12968));
    defparam i10861_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i10881_3_lut (.I0(rd_addr_p1cmp_r[2]), .I1(n12968), .I2(wr_addr_r[2]), 
            .I3(GND_net), .O(n12990));
    defparam i10881_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 i10936_4_lut (.I0(\MISC.wr_w ), .I1(n12990), .I2(rd_addr_p1cmp_r[3]), 
            .I3(wr_addr_r[3]), .O(n13046));
    defparam i10936_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i2_3_lut_adj_62 (.I0(\MISC.empty_flag_r ), .I1(DEBUG_2_c), .I2(full_nxt_w_N_812), 
            .I3(GND_net), .O(empty_nxt_w_N_823));
    defparam i2_3_lut_adj_62.LUT_INIT = 16'h0202;
    SB_LUT4 i5250_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[6] ), 
            .I3(\mem_REG.mem_3_6 ), .O(n6724));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5250_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15475_bdd_4_lut (.I0(n15475), .I1(n13700), .I2(n13699), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[23]));
    defparam n15475_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14587_bdd_4_lut (.I0(n14587), .I1(\mem_REG.mem_1_4 ), .I2(\mem_REG.mem_0_4 ), 
            .I3(rd_addr_r[1]), .O(n14590));
    defparam n14587_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5249_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[5] ), 
            .I3(\mem_REG.mem_3_5 ), .O(n6723));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5249_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_63 (.I0(reset_all), .I1(\MISC.rd_w ), .I2(empty_nxt_w_N_823), 
            .I3(n13046), .O(empty_ext_r_N_796));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i1_4_lut_adj_63.LUT_INIT = 16'hfafe;
    SB_LUT4 i5248_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[4] ), 
            .I3(\mem_REG.mem_3_4 ), .O(n6722));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5248_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_64 (.I0(wr_addr_r[2]), .I1(\MISC.wr_flag_addr_r [0]), 
            .I2(rd_addr_r[2]), .I3(\MISC.rd_flag_addr_r [0]), .O(n4_adj_1367));   // src/fifo_sc_32_lut_gen.v(136[186:216])
    defparam i1_4_lut_adj_64.LUT_INIT = 16'h7bde;
    SB_LUT4 i5247_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[3] ), 
            .I3(\mem_REG.mem_3_3 ), .O(n6721));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5247_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_65 (.I0(wr_addr_r[1]), .I1(n4_adj_1367), .I2(rd_addr_r[1]), 
            .I3(GND_net), .O(full_nxt_w_N_812));   // src/fifo_sc_32_lut_gen.v(136[186:216])
    defparam i2_3_lut_adj_65.LUT_INIT = 16'hdede;
    SB_LUT4 i2_4_lut_adj_66 (.I0(wr_addr_p1_r[3]), .I1(wr_cmpaddr_p1_r[1]), 
            .I2(rd_addr_r[3]), .I3(rd_addr_r[1]), .O(n6_adj_1368));
    defparam i2_4_lut_adj_66.LUT_INIT = 16'h4812;
    SB_LUT4 i10865_4_lut (.I0(\MISC.wr_flag_addr_p1_r [0]), .I1(wr_cmpaddr_p1_r[2]), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(rd_addr_r[2]), .O(n12972));
    defparam i10865_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_3_lut_adj_67 (.I0(n12972), .I1(n2057), .I2(n6_adj_1368), 
            .I3(GND_net), .O(full_nxt_w_N_797));
    defparam i2_3_lut_adj_67.LUT_INIT = 16'h4040;
    SB_LUT4 i7221_4_lut (.I0(full_nxt_w_N_797), .I1(reset_all), .I2(\MISC.full_flag_r ), 
            .I3(n12934), .O(full_ext_r_N_794));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7221_4_lut.LUT_INIT = 16'h2232;
    SB_LUT4 i5246_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[2] ), 
            .I3(\mem_REG.mem_3_2 ), .O(n6720));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5246_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5245_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[1] ), 
            .I3(\mem_REG.mem_3_1 ), .O(n6719));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5245_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5244_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(DEBUG_5_c_0), 
            .I3(\mem_REG.mem_3_0 ), .O(n6718));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5244_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5243_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[31] ), 
            .I3(\mem_REG.mem_2_31 ), .O(n6717));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5243_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5242_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[30] ), 
            .I3(\mem_REG.mem_2_30 ), .O(n6716));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5242_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5241_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[29] ), 
            .I3(\mem_REG.mem_2_29 ), .O(n6715));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5241_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5240_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[28] ), 
            .I3(\mem_REG.mem_2_28 ), .O(n6714));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5240_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5239_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[27] ), 
            .I3(\mem_REG.mem_2_27 ), .O(n6713));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5239_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7226_2_lut (.I0(rd_addr_nxt_w[0]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(rd_addr_p1_r_3__N_712[0]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7226_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i5238_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[26] ), 
            .I3(\mem_REG.mem_2_26 ), .O(n6712));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5238_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5237_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[25] ), 
            .I3(\mem_REG.mem_2_25 ), .O(n6711));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5237_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5236_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[24] ), 
            .I3(\mem_REG.mem_2_24 ), .O(n6710));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5236_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \mem_REG.data_raw_r_i0_i2  (.Q(sc32_fifo_data_out[1]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[1]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_LUT4 i5235_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[23] ), 
            .I3(\mem_REG.mem_2_23 ), .O(n6709));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5235_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5234_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[22] ), 
            .I3(\mem_REG.mem_2_22 ), .O(n6708));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5234_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5233_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[21] ), 
            .I3(\mem_REG.mem_2_21 ), .O(n6707));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5233_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_12902  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_12 ), .I2(\mem_REG.mem_3_12 ), .I3(rd_addr_r[1]), 
            .O(n14737));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_12902 .LUT_INIT = 16'he4aa;
    SB_LUT4 n14737_bdd_4_lut (.I0(n14737), .I1(\mem_REG.mem_1_12 ), .I2(\mem_REG.mem_0_12 ), 
            .I3(rd_addr_r[1]), .O(n14740));
    defparam n14737_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12722 (.I0(rd_addr_r[1]), .I1(n13132), 
            .I2(n13133), .I3(rd_addr_r[2]), .O(n14731));
    defparam rd_addr_r_1__bdd_4_lut_12722.LUT_INIT = 16'he4aa;
    SB_LUT4 n14731_bdd_4_lut (.I0(n14731), .I1(n13130), .I2(n13129), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[0]));
    defparam n14731_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13196 (.I0(rd_addr_r[1]), .I1(n13663), 
            .I2(n13664), .I3(rd_addr_r[2]), .O(n15451));
    defparam rd_addr_r_1__bdd_4_lut_13196.LUT_INIT = 16'he4aa;
    SB_LUT4 n15451_bdd_4_lut (.I0(n15451), .I1(n13646), .I2(n13645), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[21]));
    defparam n15451_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7225_2_lut (.I0(rd_addr_nxt_w[0]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(rd_addr_r_3__N_708[0]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7225_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5232_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[20] ), 
            .I3(\mem_REG.mem_2_20 ), .O(n6706));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5232_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7223_2_lut (.I0(wr_addr_nxt_w[0]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(wr_addr_p1_r_3__N_694[0]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7223_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i5231_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[19] ), 
            .I3(\mem_REG.mem_2_19 ), .O(n6705));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5231_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5230_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[18] ), 
            .I3(\mem_REG.mem_2_18 ), .O(n6704));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5230_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_en_i_I_0_180_2_lut (.I0(DEBUG_2_c), .I1(\MISC.full_flag_r ), 
            .I2(GND_net), .I3(GND_net), .O(\MISC.wr_w ));   // src/fifo_sc_32_lut_gen.v(268[25:51])
    defparam wr_en_i_I_0_180_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5229_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[17] ), 
            .I3(\mem_REG.mem_2_17 ), .O(n6703));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5229_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13176 (.I0(rd_addr_r[1]), .I1(n13813), 
            .I2(n13814), .I3(rd_addr_r[2]), .O(n15433));
    defparam rd_addr_r_1__bdd_4_lut_13176.LUT_INIT = 16'he4aa;
    SB_LUT4 n15433_bdd_4_lut (.I0(n15433), .I1(n13637), .I2(n13636), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[7]));
    defparam n15433_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5228_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[16] ), 
            .I3(\mem_REG.mem_2_16 ), .O(n6702));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5228_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5227_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[15] ), 
            .I3(\mem_REG.mem_2_15 ), .O(n6701));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5227_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5226_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[14] ), 
            .I3(\mem_REG.mem_2_14 ), .O(n6700));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5226_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5225_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[13] ), 
            .I3(\mem_REG.mem_2_13 ), .O(n6699));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5225_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7218_2_lut (.I0(wr_addr_nxt_w[0]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(wr_addr_r_3__N_690[0]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7218_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE \mem_REG.data_raw_r_i0_i3  (.Q(sc32_fifo_data_out[2]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[2]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_LUT4 i5224_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[12] ), 
            .I3(\mem_REG.mem_2_12 ), .O(n6698));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5224_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5223_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[11] ), 
            .I3(\mem_REG.mem_2_11 ), .O(n6697));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5223_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5222_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[10] ), 
            .I3(\mem_REG.mem_2_10 ), .O(n6696));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5222_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5221_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[9] ), 
            .I3(\mem_REG.mem_2_9 ), .O(n6695));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5221_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5220_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[8] ), 
            .I3(\mem_REG.mem_2_8 ), .O(n6694));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5220_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5219_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[7] ), 
            .I3(\mem_REG.mem_2_7 ), .O(n6693));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5219_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11672_3_lut (.I0(\mem_REG.mem_0_27 ), .I1(\mem_REG.mem_1_27 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13783));
    defparam i11672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11673_3_lut (.I0(\mem_REG.mem_2_27 ), .I1(\mem_REG.mem_3_27 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13784));
    defparam i11673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5218_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[6] ), 
            .I3(\mem_REG.mem_2_6 ), .O(n6692));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5218_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5217_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[5] ), 
            .I3(\mem_REG.mem_2_5 ), .O(n6691));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5217_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11697_3_lut (.I0(\mem_REG.mem_6_27 ), .I1(\mem_REG.mem_7_27 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13808));
    defparam i11697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5216_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[4] ), 
            .I3(\mem_REG.mem_2_4 ), .O(n6690));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5216_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11696_3_lut (.I0(\mem_REG.mem_4_27 ), .I1(\mem_REG.mem_5_27 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13807));
    defparam i11696_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE \mem_REG.data_raw_r_i0_i4  (.Q(sc32_fifo_data_out[3]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[3]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i5  (.Q(sc32_fifo_data_out[4]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[4]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i6  (.Q(sc32_fifo_data_out[5]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[5]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i7  (.Q(sc32_fifo_data_out[6]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[6]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i8  (.Q(sc32_fifo_data_out[7]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[7]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i9  (.Q(sc32_fifo_data_out[8]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[8]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i10  (.Q(sc32_fifo_data_out[9]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[9]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i11  (.Q(sc32_fifo_data_out[10]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[10]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i12  (.Q(sc32_fifo_data_out[11]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[11]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i13  (.Q(sc32_fifo_data_out[12]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[12]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i14  (.Q(sc32_fifo_data_out[13]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[13]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i15  (.Q(sc32_fifo_data_out[14]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[14]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i16  (.Q(sc32_fifo_data_out[15]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[15]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i17  (.Q(sc32_fifo_data_out[16]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[16]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i18  (.Q(sc32_fifo_data_out[17]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[17]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i19  (.Q(sc32_fifo_data_out[18]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[18]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i20  (.Q(sc32_fifo_data_out[19]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[19]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i21  (.Q(sc32_fifo_data_out[20]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[20]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i22  (.Q(sc32_fifo_data_out[21]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[21]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i23  (.Q(sc32_fifo_data_out[22]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[22]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i24  (.Q(sc32_fifo_data_out[23]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[23]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i25  (.Q(sc32_fifo_data_out[24]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[24]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i26  (.Q(sc32_fifo_data_out[25]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[25]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i27  (.Q(sc32_fifo_data_out[26]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[26]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i28  (.Q(sc32_fifo_data_out[27]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[27]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i29  (.Q(sc32_fifo_data_out[28]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[28]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i30  (.Q(sc32_fifo_data_out[29]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[29]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i31  (.Q(sc32_fifo_data_out[30]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[30]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i32  (.Q(sc32_fifo_data_out[31]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[31]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13161 (.I0(rd_addr_r[1]), .I1(n13702), 
            .I2(n13703), .I3(rd_addr_r[2]), .O(n15409));
    defparam rd_addr_r_1__bdd_4_lut_13161.LUT_INIT = 16'he4aa;
    SB_LUT4 n15409_bdd_4_lut (.I0(n15409), .I1(n13622), .I2(n13621), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[20]));
    defparam n15409_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_14 ), .I2(\mem_REG.mem_3_14 ), .I3(rd_addr_r[1]), 
            .O(n16201));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut .LUT_INIT = 16'he4aa;
    SB_LUT4 i5215_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[3] ), 
            .I3(\mem_REG.mem_2_3 ), .O(n6689));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5215_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5214_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[2] ), 
            .I3(\mem_REG.mem_2_2 ), .O(n6688));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5214_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5213_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[1] ), 
            .I3(\mem_REG.mem_2_1 ), .O(n6687));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5213_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11669_3_lut (.I0(\mem_REG.mem_0_10 ), .I1(\mem_REG.mem_1_10 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13780));
    defparam i11669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11670_3_lut (.I0(\mem_REG.mem_2_10 ), .I1(\mem_REG.mem_3_10 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13781));
    defparam i11670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5212_3_lut_4_lut (.I0(n6), .I1(wr_addr_r[2]), .I2(DEBUG_5_c_0), 
            .I3(\mem_REG.mem_2_0 ), .O(n6686));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5212_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16201_bdd_4_lut (.I0(n16201), .I1(\mem_REG.mem_1_14 ), .I2(\mem_REG.mem_0_14 ), 
            .I3(rd_addr_r[1]), .O(n16204));
    defparam n16201_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11691_3_lut (.I0(\mem_REG.mem_6_10 ), .I1(\mem_REG.mem_7_10 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13802));
    defparam i11691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5211_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[31] ), 
            .I3(\mem_REG.mem_1_31 ), .O(n6685));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5211_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5210_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[30] ), 
            .I3(\mem_REG.mem_1_30 ), .O(n6684));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5210_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11690_3_lut (.I0(\mem_REG.mem_4_10 ), .I1(\mem_REG.mem_5_10 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13801));
    defparam i11690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5209_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[29] ), 
            .I3(\mem_REG.mem_1_29 ), .O(n6683));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5209_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5208_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[28] ), 
            .I3(\mem_REG.mem_1_28 ), .O(n6682));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5208_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5207_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[27] ), 
            .I3(\mem_REG.mem_1_27 ), .O(n6681));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5207_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5206_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[26] ), 
            .I3(\mem_REG.mem_1_26 ), .O(n6680));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5206_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5205_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[25] ), 
            .I3(\mem_REG.mem_1_25 ), .O(n6679));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5205_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5204_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[24] ), 
            .I3(\mem_REG.mem_1_24 ), .O(n6678));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5204_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF wr_addr_r_i1 (.Q(wr_addr_r[1]), .C(SLM_CLK_c), .D(wr_addr_r_3__N_690[1]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_LUT4 i5203_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[23] ), 
            .I3(\mem_REG.mem_1_23 ), .O(n6677));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5203_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5202_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[22] ), 
            .I3(\mem_REG.mem_1_22 ), .O(n6676));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5202_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5201_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[21] ), 
            .I3(\mem_REG.mem_1_21 ), .O(n6675));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5201_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5200_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[20] ), 
            .I3(\mem_REG.mem_1_20 ), .O(n6674));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5200_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF wr_addr_r_i2 (.Q(wr_addr_r[2]), .C(SLM_CLK_c), .D(wr_addr_r_3__N_690[2]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_LUT4 i5199_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[19] ), 
            .I3(\mem_REG.mem_1_19 ), .O(n6673));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5199_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5198_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[18] ), 
            .I3(\mem_REG.mem_1_18 ), .O(n6672));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5198_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5197_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[17] ), 
            .I3(\mem_REG.mem_1_17 ), .O(n6671));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5197_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF wr_addr_r_i3 (.Q(wr_addr_r[3]), .C(SLM_CLK_c), .D(wr_addr_r_3__N_690[3]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF wr_addr_p1_r_i3 (.Q(wr_addr_p1_r[3]), .C(SLM_CLK_c), .D(wr_addr_p1cmp_r_3__N_698[3]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF wr_cmpaddr_p1_r_i1 (.Q(wr_cmpaddr_p1_r[1]), .C(SLM_CLK_c), .D(wr_addr_p1_r_3__N_694[1]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF wr_cmpaddr_p1_r_i2 (.Q(wr_cmpaddr_p1_r[2]), .C(SLM_CLK_c), .D(wr_addr_p1_r_3__N_694[2]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF rd_addr_r_i1 (.Q(rd_addr_r[1]), .C(SLM_CLK_c), .D(rd_addr_r_3__N_708[1]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF rd_addr_r_i2 (.Q(rd_addr_r[2]), .C(SLM_CLK_c), .D(rd_addr_r_3__N_708[2]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF rd_addr_r_i3 (.Q(rd_addr_r[3]), .C(SLM_CLK_c), .D(rd_addr_r_3__N_708[3]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF rd_addr_p1cmp_r_i1 (.Q(rd_addr_p1cmp_r[1]), .C(SLM_CLK_c), .D(rd_addr_p1_r_3__N_712[1]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF rd_addr_p1cmp_r_i2 (.Q(rd_addr_p1cmp_r[2]), .C(SLM_CLK_c), .D(rd_addr_p1_r_3__N_712[2]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF rd_addr_p1cmp_r_i3 (.Q(rd_addr_p1cmp_r[3]), .C(SLM_CLK_c), .D(rd_addr_p1_r_3__N_712[3]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_LUT4 i5196_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[16] ), 
            .I3(\mem_REG.mem_1_16 ), .O(n6670));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5196_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5195_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[15] ), 
            .I3(\mem_REG.mem_1_15 ), .O(n6669));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5195_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5194_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[14] ), 
            .I3(\mem_REG.mem_1_14 ), .O(n6668));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5194_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5193_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[13] ), 
            .I3(\mem_REG.mem_1_13 ), .O(n6667));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5193_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5192_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[12] ), 
            .I3(\mem_REG.mem_1_12 ), .O(n6666));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5192_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5191_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[11] ), 
            .I3(\mem_REG.mem_1_11 ), .O(n6665));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5191_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5190_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[10] ), 
            .I3(\mem_REG.mem_1_10 ), .O(n6664));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5190_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5189_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[9] ), 
            .I3(\mem_REG.mem_1_9 ), .O(n6663));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5189_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5188_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[8] ), 
            .I3(\mem_REG.mem_1_8 ), .O(n6662));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5188_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_13800  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_15 ), .I2(\mem_REG.mem_7_15 ), .I3(rd_addr_r[1]), 
            .O(n16159));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_13800 .LUT_INIT = 16'he4aa;
    SB_LUT4 i5187_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[7] ), 
            .I3(\mem_REG.mem_1_7 ), .O(n6661));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5187_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5186_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[6] ), 
            .I3(\mem_REG.mem_1_6 ), .O(n6660));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5186_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16159_bdd_4_lut (.I0(n16159), .I1(\mem_REG.mem_5_15 ), .I2(\mem_REG.mem_4_15 ), 
            .I3(rd_addr_r[1]), .O(n16162));
    defparam n16159_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13141 (.I0(rd_addr_r[1]), .I1(n13816), 
            .I2(n13817), .I3(rd_addr_r[2]), .O(n15373));
    defparam rd_addr_r_1__bdd_4_lut_13141.LUT_INIT = 16'he4aa;
    SB_LUT4 i5185_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[5] ), 
            .I3(\mem_REG.mem_1_5 ), .O(n6659));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5185_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5184_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[4] ), 
            .I3(\mem_REG.mem_1_4 ), .O(n6658));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5184_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15373_bdd_4_lut (.I0(n15373), .I1(n13574), .I2(n13573), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[6]));
    defparam n15373_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5183_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[3] ), 
            .I3(\mem_REG.mem_1_3 ), .O(n6657));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5183_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5182_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[2] ), 
            .I3(\mem_REG.mem_1_2 ), .O(n6656));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5182_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5181_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[1] ), 
            .I3(\mem_REG.mem_1_1 ), .O(n6655));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5181_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5180_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(DEBUG_5_c_0), 
            .I3(\mem_REG.mem_1_0 ), .O(n6654));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5180_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5179_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[31] ), 
            .I3(\mem_REG.mem_0_31 ), .O(n6653));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5179_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5178_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[30] ), 
            .I3(\mem_REG.mem_0_30 ), .O(n6652));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5178_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5177_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[29] ), 
            .I3(\mem_REG.mem_0_29 ), .O(n6651));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5177_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5176_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[28] ), 
            .I3(\mem_REG.mem_0_28 ), .O(n6650));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5176_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5175_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[27] ), 
            .I3(\mem_REG.mem_0_27 ), .O(n6649));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5175_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5174_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[26] ), 
            .I3(\mem_REG.mem_0_26 ), .O(n6648));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5174_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_13765  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_31 ), .I2(\mem_REG.mem_7_31 ), .I3(rd_addr_r[1]), 
            .O(n16063));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_13765 .LUT_INIT = 16'he4aa;
    SB_LUT4 n16063_bdd_4_lut (.I0(n16063), .I1(\mem_REG.mem_5_31 ), .I2(\mem_REG.mem_4_31 ), 
            .I3(rd_addr_r[1]), .O(n16066));
    defparam n16063_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5173_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[25] ), 
            .I3(\mem_REG.mem_0_25 ), .O(n6647));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5173_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5172_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[24] ), 
            .I3(\mem_REG.mem_0_24 ), .O(n6646));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5172_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5171_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[23] ), 
            .I3(\mem_REG.mem_0_23 ), .O(n6645));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5171_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5170_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[22] ), 
            .I3(\mem_REG.mem_0_22 ), .O(n6644));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5170_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5169_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[21] ), 
            .I3(\mem_REG.mem_0_21 ), .O(n6643));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5169_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5168_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[20] ), 
            .I3(\mem_REG.mem_0_20 ), .O(n6642));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5168_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5167_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[19] ), 
            .I3(\mem_REG.mem_0_19 ), .O(n6641));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5167_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5166_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[18] ), 
            .I3(\mem_REG.mem_0_18 ), .O(n6640));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5166_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5165_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[17] ), 
            .I3(\mem_REG.mem_0_17 ), .O(n6639));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5165_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5164_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[16] ), 
            .I3(\mem_REG.mem_0_16 ), .O(n6638));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5164_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_en_i_I_0_181_2_lut (.I0(sc32_fifo_read_enable), .I1(\MISC.empty_flag_r ), 
            .I2(GND_net), .I3(GND_net), .O(\MISC.rd_w ));   // src/fifo_sc_32_lut_gen.v(269[25:52])
    defparam rd_en_i_I_0_181_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5163_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[15] ), 
            .I3(\mem_REG.mem_0_15 ), .O(n6637));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5163_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5162_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[14] ), 
            .I3(\mem_REG.mem_0_14 ), .O(n6636));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5162_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5161_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[13] ), 
            .I3(\mem_REG.mem_0_13 ), .O(n6635));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5161_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5160_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[12] ), 
            .I3(\mem_REG.mem_0_12 ), .O(n6634));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5160_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5159_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[11] ), 
            .I3(\mem_REG.mem_0_11 ), .O(n6633));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5159_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5158_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[10] ), 
            .I3(\mem_REG.mem_0_10 ), .O(n6632));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5158_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_13366  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_30 ), .I2(\mem_REG.mem_3_30 ), .I3(rd_addr_r[1]), 
            .O(n15283));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_13366 .LUT_INIT = 16'he4aa;
    SB_LUT4 i5157_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[9] ), 
            .I3(\mem_REG.mem_0_9 ), .O(n6631));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5157_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5156_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[8] ), 
            .I3(\mem_REG.mem_0_8 ), .O(n6630));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5156_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5155_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[7] ), 
            .I3(\mem_REG.mem_0_7 ), .O(n6629));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5155_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5154_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[6] ), 
            .I3(\mem_REG.mem_0_6 ), .O(n6628));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5154_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5153_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[5] ), 
            .I3(\mem_REG.mem_0_5 ), .O(n6627));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5153_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15283_bdd_4_lut (.I0(n15283), .I1(\mem_REG.mem_1_30 ), .I2(\mem_REG.mem_0_30 ), 
            .I3(rd_addr_r[1]), .O(n15286));
    defparam n15283_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_13036  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_30 ), .I2(\mem_REG.mem_7_30 ), .I3(rd_addr_r[1]), 
            .O(n15259));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_13036 .LUT_INIT = 16'he4aa;
    SB_LUT4 n15259_bdd_4_lut (.I0(n15259), .I1(\mem_REG.mem_5_30 ), .I2(\mem_REG.mem_4_30 ), 
            .I3(rd_addr_r[1]), .O(n15262));
    defparam n15259_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5152_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[4] ), 
            .I3(\mem_REG.mem_0_4 ), .O(n6626));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5152_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5151_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[3] ), 
            .I3(\mem_REG.mem_0_3 ), .O(n6625));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5151_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5150_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[2] ), 
            .I3(\mem_REG.mem_0_2 ), .O(n6624));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5150_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5149_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(\dc32_fifo_data_out[1] ), 
            .I3(\mem_REG.mem_0_1 ), .O(n6623));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5149_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5148_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(DEBUG_5_c_0), 
            .I3(\mem_REG.mem_0_0 ), .O(n6622));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5148_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_13685  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_29 ), .I2(\mem_REG.mem_7_29 ), .I3(rd_addr_r[1]), 
            .O(n15985));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_13685 .LUT_INIT = 16'he4aa;
    SB_LUT4 n15985_bdd_4_lut (.I0(n15985), .I1(\mem_REG.mem_5_29 ), .I2(\mem_REG.mem_4_29 ), 
            .I3(rd_addr_r[1]), .O(n15988));
    defparam n15985_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_13016  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_31 ), .I2(\mem_REG.mem_3_31 ), .I3(rd_addr_r[1]), 
            .O(n15211));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_13016 .LUT_INIT = 16'he4aa;
    SB_LUT4 n15211_bdd_4_lut (.I0(n15211), .I1(\mem_REG.mem_1_31 ), .I2(\mem_REG.mem_0_31 ), 
            .I3(rd_addr_r[1]), .O(n15214));
    defparam n15211_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_12976  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_5 ), .I2(\mem_REG.mem_3_5 ), .I3(rd_addr_r[1]), 
            .O(n15193));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_12976 .LUT_INIT = 16'he4aa;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_12458  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_5 ), .I2(\mem_REG.mem_7_5 ), .I3(rd_addr_r[1]), 
            .O(n14569));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_12458 .LUT_INIT = 16'he4aa;
    SB_LUT4 n15193_bdd_4_lut (.I0(n15193), .I1(\mem_REG.mem_1_5 ), .I2(\mem_REG.mem_0_5 ), 
            .I3(rd_addr_r[1]), .O(n15196));
    defparam n15193_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut (.I0(rd_addr_r[1]), .I1(n14203), .I2(n14204), 
            .I3(rd_addr_r[2]), .O(n15925));
    defparam rd_addr_r_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n15925_bdd_4_lut (.I0(n15925), .I1(n14192), .I2(n14191), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[17]));
    defparam n15925_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13571 (.I0(rd_addr_r[1]), .I1(n14185), 
            .I2(n14186), .I3(rd_addr_r[2]), .O(n15919));
    defparam rd_addr_r_1__bdd_4_lut_13571.LUT_INIT = 16'he4aa;
    SB_LUT4 n15919_bdd_4_lut (.I0(n15919), .I1(n14168), .I2(n14167), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[16]));
    defparam n15919_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14569_bdd_4_lut (.I0(n14569), .I1(\mem_REG.mem_5_5 ), .I2(\mem_REG.mem_4_5 ), 
            .I3(rd_addr_r[1]), .O(n14572));
    defparam n14569_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_12961  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_1 ), .I2(\mem_REG.mem_3_1 ), .I3(rd_addr_r[1]), 
            .O(n15121));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_12961 .LUT_INIT = 16'he4aa;
    SB_LUT4 n15121_bdd_4_lut (.I0(n15121), .I1(\mem_REG.mem_1_1 ), .I2(\mem_REG.mem_0_1 ), 
            .I3(rd_addr_r[1]), .O(n15124));
    defparam n15121_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_13621  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_15 ), .I2(\mem_REG.mem_3_15 ), .I3(rd_addr_r[1]), 
            .O(n15853));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_13621 .LUT_INIT = 16'he4aa;
    SB_LUT4 n15853_bdd_4_lut (.I0(n15853), .I1(\mem_REG.mem_1_15 ), .I2(\mem_REG.mem_0_15 ), 
            .I3(rd_addr_r[1]), .O(n15856));
    defparam n15853_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_13511  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_14 ), .I2(\mem_REG.mem_7_14 ), .I3(rd_addr_r[1]), 
            .O(n15835));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_13511 .LUT_INIT = 16'he4aa;
    SB_LUT4 n15835_bdd_4_lut (.I0(n15835), .I1(\mem_REG.mem_5_14 ), .I2(\mem_REG.mem_4_14 ), 
            .I3(rd_addr_r[1]), .O(n15838));
    defparam n15835_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_13496  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_12 ), .I2(\mem_REG.mem_7_12 ), .I3(rd_addr_r[1]), 
            .O(n15811));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_13496 .LUT_INIT = 16'he4aa;
    SB_LUT4 n15811_bdd_4_lut (.I0(n15811), .I1(\mem_REG.mem_5_12 ), .I2(\mem_REG.mem_4_12 ), 
            .I3(rd_addr_r[1]), .O(n15814));
    defparam n15811_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_13111 (.I0(rd_addr_r[1]), .I1(n13456), 
            .I2(n13457), .I3(rd_addr_r[2]), .O(n15079));
    defparam rd_addr_r_1__bdd_4_lut_13111.LUT_INIT = 16'he4aa;
    SB_LUT4 n15079_bdd_4_lut (.I0(n15079), .I1(n13334), .I2(n13333), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[3]));
    defparam n15079_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_13476  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_11 ), .I2(\mem_REG.mem_7_11 ), .I3(rd_addr_r[1]), 
            .O(n15799));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_13476 .LUT_INIT = 16'he4aa;
    SB_LUT4 n15799_bdd_4_lut (.I0(n15799), .I1(\mem_REG.mem_5_11 ), .I2(\mem_REG.mem_4_11 ), 
            .I3(rd_addr_r[1]), .O(n15802));
    defparam n15799_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11576_3_lut (.I0(\mem_REG.mem_4_22 ), .I1(\mem_REG.mem_5_22 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13687));
    defparam i11576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11577_3_lut (.I0(\mem_REG.mem_6_22 ), .I1(\mem_REG.mem_7_22 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13688));
    defparam i11577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11565_3_lut (.I0(\mem_REG.mem_2_22 ), .I1(\mem_REG.mem_3_22 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13676));
    defparam i11565_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11564_3_lut (.I0(\mem_REG.mem_0_22 ), .I1(\mem_REG.mem_1_22 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13675));
    defparam i11564_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7384_3_lut_4_lut (.I0(rd_addr_nxt_w[2]), .I1(reset_all), .I2(rd_addr_nxt_w[1]), 
            .I3(rd_addr_nxt_w[0]), .O(rd_addr_p1_r_3__N_712[2]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7384_3_lut_4_lut.LUT_INIT = 16'h1222;
    SB_LUT4 rd_addr_r_3__I_0_i4_3_lut_4_lut (.I0(rd_addr_r[3]), .I1(rd_addr_p1cmp_r[3]), 
            .I2(sc32_fifo_read_enable), .I3(\MISC.empty_flag_r ), .O(rd_addr_nxt_w[3]));   // src/fifo_sc_32_lut_gen.v(133[44:95])
    defparam rd_addr_r_3__I_0_i4_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7382_2_lut_4_lut (.I0(rd_addr_r[3]), .I1(rd_addr_p1cmp_r[3]), 
            .I2(\MISC.rd_w ), .I3(reset_all), .O(rd_addr_r_3__N_708[3]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7382_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 rd_addr_r_3__I_0_i3_3_lut_4_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1cmp_r[2]), 
            .I2(sc32_fifo_read_enable), .I3(\MISC.empty_flag_r ), .O(rd_addr_nxt_w[2]));   // src/fifo_sc_32_lut_gen.v(133[44:95])
    defparam rd_addr_r_3__I_0_i3_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 rd_addr_r_3__I_0_i2_3_lut_4_lut (.I0(rd_addr_r[1]), .I1(rd_addr_p1cmp_r[1]), 
            .I2(sc32_fifo_read_enable), .I3(\MISC.empty_flag_r ), .O(rd_addr_nxt_w[1]));   // src/fifo_sc_32_lut_gen.v(133[44:95])
    defparam rd_addr_r_3__I_0_i2_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7379_3_lut_4_lut (.I0(wr_addr_nxt_w[2]), .I1(reset_all), .I2(wr_addr_nxt_w[1]), 
            .I3(wr_addr_nxt_w[0]), .O(wr_addr_p1_r_3__N_694[2]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7379_3_lut_4_lut.LUT_INIT = 16'h1222;
    SB_LUT4 wr_addr_r_3__I_0_i4_3_lut_4_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_r[3]), 
            .I2(DEBUG_2_c), .I3(\MISC.full_flag_r ), .O(wr_addr_nxt_w[3]));   // src/fifo_sc_32_lut_gen.v(130[44:94])
    defparam wr_addr_r_3__I_0_i4_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7377_2_lut_4_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_r[3]), 
            .I2(\MISC.wr_w ), .I3(reset_all), .O(wr_addr_r_3__N_690[3]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7377_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 i11603_3_lut (.I0(\mem_REG.mem_4_23 ), .I1(\mem_REG.mem_5_23 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13714));
    defparam i11603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11604_3_lut (.I0(\mem_REG.mem_6_23 ), .I1(\mem_REG.mem_7_23 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13715));
    defparam i11604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_3__I_0_i3_3_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_cmpaddr_p1_r[2]), 
            .I2(DEBUG_2_c), .I3(\MISC.full_flag_r ), .O(wr_addr_nxt_w[2]));   // src/fifo_sc_32_lut_gen.v(130[44:94])
    defparam wr_addr_r_3__I_0_i3_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 wr_addr_r_3__I_0_i2_3_lut_4_lut (.I0(wr_addr_r[1]), .I1(wr_cmpaddr_p1_r[1]), 
            .I2(DEBUG_2_c), .I3(\MISC.full_flag_r ), .O(wr_addr_nxt_w[1]));   // src/fifo_sc_32_lut_gen.v(130[44:94])
    defparam wr_addr_r_3__I_0_i2_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i2218_3_lut_4_lut_4_lut (.I0(DEBUG_2_c), .I1(\MISC.full_flag_r ), 
            .I2(sc32_fifo_read_enable), .I3(\MISC.empty_flag_r ), .O(n3679));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i2218_3_lut_4_lut_4_lut.LUT_INIT = 16'h00d0;
    SB_LUT4 i11589_3_lut (.I0(\mem_REG.mem_2_23 ), .I1(\mem_REG.mem_3_23 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13700));
    defparam i11589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11588_3_lut (.I0(\mem_REG.mem_0_23 ), .I1(\mem_REG.mem_1_23 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13699));
    defparam i11588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7739115_i1_3_lut (.I0(n15124), .I1(n15700), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[1]));
    defparam i7739115_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11021_3_lut (.I0(\mem_REG.mem_4_0 ), .I1(\mem_REG.mem_5_0 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13132));
    defparam i11021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11022_3_lut (.I0(\mem_REG.mem_6_0 ), .I1(\mem_REG.mem_7_0 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13133));
    defparam i11022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11019_3_lut (.I0(\mem_REG.mem_2_0 ), .I1(\mem_REG.mem_3_0 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13130));
    defparam i11019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11018_3_lut (.I0(\mem_REG.mem_0_0 ), .I1(\mem_REG.mem_1_0 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13129));
    defparam i11018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11552_3_lut (.I0(\mem_REG.mem_4_21 ), .I1(\mem_REG.mem_5_21 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13663));
    defparam i11552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11553_3_lut (.I0(\mem_REG.mem_6_21 ), .I1(\mem_REG.mem_7_21 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13664));
    defparam i11553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11535_3_lut (.I0(\mem_REG.mem_2_21 ), .I1(\mem_REG.mem_3_21 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13646));
    defparam i11535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11534_3_lut (.I0(\mem_REG.mem_0_21 ), .I1(\mem_REG.mem_1_21 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13645));
    defparam i11534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11702_3_lut (.I0(\mem_REG.mem_4_7 ), .I1(\mem_REG.mem_5_7 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13813));
    defparam i11702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11703_3_lut (.I0(\mem_REG.mem_6_7 ), .I1(\mem_REG.mem_7_7 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13814));
    defparam i11703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11526_3_lut (.I0(\mem_REG.mem_2_7 ), .I1(\mem_REG.mem_3_7 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13637));
    defparam i11526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11525_3_lut (.I0(\mem_REG.mem_0_7 ), .I1(\mem_REG.mem_1_7 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13636));
    defparam i11525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7757124_i1_3_lut (.I0(n14590), .I1(n14512), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[4]));
    defparam i7757124_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7763127_i1_3_lut (.I0(n15196), .I1(n14572), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[5]));
    defparam i7763127_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7799145_i1_3_lut (.I0(n15706), .I1(n15802), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[11]));
    defparam i7799145_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7829160_i1_3_lut (.I0(n14740), .I1(n15814), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[12]));
    defparam i7829160_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7835163_i1_3_lut (.I0(n14638), .I1(n14608), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[13]));
    defparam i7835163_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7841166_i1_3_lut (.I0(n16204), .I1(n15838), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[14]));
    defparam i7841166_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7847169_i1_3_lut (.I0(n15856), .I1(n16162), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[15]));
    defparam i7847169_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7949220_i1_3_lut (.I0(n15784), .I1(n15742), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[28]));
    defparam i7949220_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7955223_i1_3_lut (.I0(n15682), .I1(n15988), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[29]));
    defparam i7955223_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7985238_i1_3_lut (.I0(n15286), .I1(n15262), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[30]));
    defparam i7985238_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7991241_i1_3_lut (.I0(n15214), .I1(n16066), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[31]));
    defparam i7991241_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11591_3_lut (.I0(\mem_REG.mem_4_20 ), .I1(\mem_REG.mem_5_20 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13702));
    defparam i11591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11592_3_lut (.I0(\mem_REG.mem_6_20 ), .I1(\mem_REG.mem_7_20 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13703));
    defparam i11592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_3__I_0_i1_3_lut_4_lut (.I0(\MISC.wr_flag_addr_r [0]), 
            .I1(\MISC.wr_flag_addr_p1_r [0]), .I2(DEBUG_2_c), .I3(\MISC.full_flag_r ), 
            .O(wr_addr_nxt_w[0]));   // src/fifo_sc_32_lut_gen.v(130[44:94])
    defparam wr_addr_r_3__I_0_i1_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 rd_addr_r_3__I_0_i1_3_lut_4_lut (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\MISC.rd_flag_addr_p1_r [0]), .I2(sc32_fifo_read_enable), 
            .I3(\MISC.empty_flag_r ), .O(rd_addr_nxt_w[0]));   // src/fifo_sc_32_lut_gen.v(133[44:95])
    defparam rd_addr_r_3__I_0_i1_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i11511_3_lut (.I0(\mem_REG.mem_2_20 ), .I1(\mem_REG.mem_3_20 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13622));
    defparam i11511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11510_3_lut (.I0(\mem_REG.mem_0_20 ), .I1(\mem_REG.mem_1_20 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13621));
    defparam i11510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10827_2_lut_4_lut (.I0(sc32_fifo_read_enable), .I1(wr_addr_r[1]), 
            .I2(n4_adj_1367), .I3(rd_addr_r[1]), .O(n12934));
    defparam i10827_2_lut_4_lut.LUT_INIT = 16'hfbfe;
    SB_LUT4 i1036_2_lut_4_lut (.I0(sc32_fifo_read_enable), .I1(\MISC.empty_flag_r ), 
            .I2(DEBUG_2_c), .I3(\MISC.full_flag_r ), .O(n2057));   // src/fifo_sc_32_lut_gen.v(270[46:60])
    defparam i1036_2_lut_4_lut.LUT_INIT = 16'h00d0;
    SB_LUT4 mux_1426_i4_3_lut_4_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_r[3]), 
            .I2(\MISC.rd_w ), .I3(\MISC.wr_w ), .O(n2775[3]));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam mux_1426_i4_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_1426_i2_3_lut_4_lut (.I0(wr_addr_r[1]), .I1(wr_cmpaddr_p1_r[1]), 
            .I2(\MISC.rd_w ), .I3(\MISC.wr_w ), .O(n2775[1]));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam mux_1426_i2_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_1426_i3_3_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_cmpaddr_p1_r[2]), 
            .I2(\MISC.rd_w ), .I3(\MISC.wr_w ), .O(n2775[2]));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam mux_1426_i3_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7375_2_lut (.I0(wr_addr_nxt_w[1]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(wr_addr_r_3__N_690[1]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7375_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7376_2_lut (.I0(wr_addr_nxt_w[2]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(wr_addr_r_3__N_690[2]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7376_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7224_4_lut (.I0(wr_addr_nxt_w[3]), .I1(reset_all), .I2(wr_addr_nxt_w[2]), 
            .I3(n3090), .O(wr_addr_p1cmp_r_3__N_698[3]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7224_4_lut.LUT_INIT = 16'h1222;
    SB_LUT4 i1646_2_lut (.I0(wr_addr_nxt_w[1]), .I1(wr_addr_nxt_w[0]), .I2(GND_net), 
            .I3(GND_net), .O(n3090));   // src/fifo_sc_32_lut_gen.v(131[47:69])
    defparam i1646_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7378_3_lut (.I0(wr_addr_nxt_w[1]), .I1(reset_all), .I2(wr_addr_nxt_w[0]), 
            .I3(GND_net), .O(wr_addr_p1_r_3__N_694[1]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7378_3_lut.LUT_INIT = 16'h1212;
    SB_LUT4 i7380_2_lut (.I0(rd_addr_nxt_w[1]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(rd_addr_r_3__N_708[1]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7380_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7381_2_lut (.I0(rd_addr_nxt_w[2]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(rd_addr_r_3__N_708[2]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7381_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7383_3_lut (.I0(rd_addr_nxt_w[1]), .I1(reset_all), .I2(rd_addr_nxt_w[0]), 
            .I3(GND_net), .O(rd_addr_p1_r_3__N_712[1]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7383_3_lut.LUT_INIT = 16'h1212;
    SB_LUT4 i1675_2_lut (.I0(rd_addr_nxt_w[1]), .I1(rd_addr_nxt_w[0]), .I2(GND_net), 
            .I3(GND_net), .O(n3119));   // src/fifo_sc_32_lut_gen.v(134[47:69])
    defparam i1675_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7385_4_lut (.I0(rd_addr_nxt_w[3]), .I1(reset_all), .I2(rd_addr_nxt_w[2]), 
            .I3(n3119), .O(rd_addr_p1_r_3__N_712[3]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i7385_4_lut.LUT_INIT = 16'h1222;
    SB_LUT4 i11705_3_lut (.I0(\mem_REG.mem_4_6 ), .I1(\mem_REG.mem_5_6 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13816));
    defparam i11705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11706_3_lut (.I0(\mem_REG.mem_6_6 ), .I1(\mem_REG.mem_7_6 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13817));
    defparam i11706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11463_3_lut (.I0(\mem_REG.mem_2_6 ), .I1(\mem_REG.mem_3_6 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13574));
    defparam i11463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11462_3_lut (.I0(\mem_REG.mem_0_6 ), .I1(\mem_REG.mem_1_6 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13573));
    defparam i11462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3893_1_lut (.I0(sc32_fifo_data_out[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5367));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3893_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3892_1_lut (.I0(sc32_fifo_data_out[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5366));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3892_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3891_1_lut (.I0(sc32_fifo_data_out[11]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5365));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3891_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3890_1_lut (.I0(sc32_fifo_data_out[12]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5364));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3890_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3889_1_lut (.I0(sc32_fifo_data_out[13]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5363));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3889_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3888_1_lut (.I0(sc32_fifo_data_out[14]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5362));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3888_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3887_1_lut (.I0(sc32_fifo_data_out[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5361));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3887_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3886_1_lut (.I0(sc32_fifo_data_out[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5360));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3886_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3885_1_lut (.I0(sc32_fifo_data_out[16]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5359));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3885_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12092_3_lut (.I0(\mem_REG.mem_4_17 ), .I1(\mem_REG.mem_5_17 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n14203));
    defparam i12092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12093_3_lut (.I0(\mem_REG.mem_6_17 ), .I1(\mem_REG.mem_7_17 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n14204));
    defparam i12093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12081_3_lut (.I0(\mem_REG.mem_2_17 ), .I1(\mem_REG.mem_3_17 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n14192));
    defparam i12081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12080_3_lut (.I0(\mem_REG.mem_0_17 ), .I1(\mem_REG.mem_1_17 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n14191));
    defparam i12080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12074_3_lut (.I0(\mem_REG.mem_4_16 ), .I1(\mem_REG.mem_5_16 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n14185));
    defparam i12074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12075_3_lut (.I0(\mem_REG.mem_6_16 ), .I1(\mem_REG.mem_7_16 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n14186));
    defparam i12075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12057_3_lut (.I0(\mem_REG.mem_2_16 ), .I1(\mem_REG.mem_3_16 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n14168));
    defparam i12057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12056_3_lut (.I0(\mem_REG.mem_0_16 ), .I1(\mem_REG.mem_1_16 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n14167));
    defparam i12056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3884_1_lut (.I0(sc32_fifo_data_out[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5358));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3884_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3883_1_lut (.I0(sc32_fifo_data_out[17]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5357));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3883_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3882_1_lut (.I0(sc32_fifo_data_out[18]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5356));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3882_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3881_1_lut (.I0(sc32_fifo_data_out[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5355));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3881_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3880_1_lut (.I0(sc32_fifo_data_out[19]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5354));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3880_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3879_1_lut (.I0(sc32_fifo_data_out[20]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5353));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3879_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3878_1_lut (.I0(sc32_fifo_data_out[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5352));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3878_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3877_1_lut (.I0(sc32_fifo_data_out[21]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5351));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3877_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3876_1_lut (.I0(sc32_fifo_data_out[22]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5350));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3876_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3875_1_lut (.I0(sc32_fifo_data_out[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5349));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3875_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3874_1_lut (.I0(sc32_fifo_data_out[23]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5348));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3874_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3873_1_lut (.I0(sc32_fifo_data_out[24]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5347));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3873_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3872_1_lut (.I0(sc32_fifo_data_out[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5346));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3872_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3871_1_lut (.I0(sc32_fifo_data_out[25]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5345));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3871_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3870_1_lut (.I0(sc32_fifo_data_out[26]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5344));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3870_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3869_1_lut (.I0(sc32_fifo_data_out[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5343));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3869_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3868_1_lut (.I0(sc32_fifo_data_out[27]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5342));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3868_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3867_1_lut (.I0(sc32_fifo_data_out[28]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5341));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3867_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3866_1_lut (.I0(sc32_fifo_data_out[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5340));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3866_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 EnabledDecoder_2_i6_2_lut_3_lut_4_lut (.I0(DEBUG_2_c), .I1(\MISC.full_flag_r ), 
            .I2(\MISC.wr_flag_addr_r [0]), .I3(wr_addr_r[1]), .O(n6));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam EnabledDecoder_2_i6_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i3865_1_lut (.I0(sc32_fifo_data_out[29]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5339));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3865_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 EnabledDecoder_2_i7_2_lut_3_lut_4_lut (.I0(DEBUG_2_c), .I1(\MISC.full_flag_r ), 
            .I2(\MISC.wr_flag_addr_r [0]), .I3(wr_addr_r[1]), .O(n7));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam EnabledDecoder_2_i7_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i3864_1_lut (.I0(sc32_fifo_data_out[30]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5338));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3864_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3863_1_lut (.I0(sc32_fifo_data_out[31]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5337));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3863_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 EnabledDecoder_2_i8_2_lut_3_lut_4_lut (.I0(DEBUG_2_c), .I1(\MISC.full_flag_r ), 
            .I2(\MISC.wr_flag_addr_r [0]), .I3(wr_addr_r[1]), .O(n8));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam EnabledDecoder_2_i8_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i9_2_lut_3_lut_4_lut (.I0(DEBUG_2_c), .I1(\MISC.full_flag_r ), 
            .I2(\MISC.wr_flag_addr_r [0]), .I3(wr_addr_r[1]), .O(n9));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam EnabledDecoder_2_i9_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i11345_3_lut (.I0(\mem_REG.mem_4_3 ), .I1(\mem_REG.mem_5_3 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13456));
    defparam i11345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11346_3_lut (.I0(\mem_REG.mem_6_3 ), .I1(\mem_REG.mem_7_3 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13457));
    defparam i11346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11223_3_lut (.I0(\mem_REG.mem_2_3 ), .I1(\mem_REG.mem_3_3 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13334));
    defparam i11223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11222_3_lut (.I0(\mem_REG.mem_0_3 ), .I1(\mem_REG.mem_1_3 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n13333));
    defparam i11222_3_lut.LUT_INIT = 16'hcaca;
>>>>>>> Stashed changes
>>>>>>> master
    
endmodule
//
// Verilog Description of module \uart_tx(CLKS_PER_BIT=20) 
//

<<<<<<< HEAD
module \uart_tx(CLKS_PER_BIT=20)  (r_SM_Main, \r_SM_Main_2__N_1025[1] , 
            UART_TX_c, SLM_CLK_c, n11691, r_Bit_Index, GND_net, n5716, 
            r_Tx_Data, n5715, n5714, n5713, \r_SM_Main_2__N_1028[0] , 
            n11079, n5712, n5711, n5710, VCC_net, n5212, n5525, 
            n5817, n5618, n5617, tx_uart_active_flag, n4715) /* synthesis syn_module_defined=1 */ ;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_1025[1] ;
=======
<<<<<<< Updated upstream
module \uart_tx(CLKS_PER_BIT=20)  (UART_TX_c, SLM_CLK_c, r_SM_Main, GND_net, 
            \r_SM_Main_2__N_841[1] , \r_SM_Main_2__N_844[0] , n3794, VCC_net, 
            n13865, n10805, n4890, r_Tx_Data, n4889, tx_uart_active_flag, 
            n5192, n5191, n5190, n5189, n5187, n5171, n5170) /* synthesis syn_module_defined=1 */ ;
>>>>>>> master
    output UART_TX_c;
    input SLM_CLK_c;
    input n11691;
    output [2:0]r_Bit_Index;
    input GND_net;
    input n5716;
    output [7:0]r_Tx_Data;
    input n5715;
    input n5714;
    input n5713;
    input \r_SM_Main_2__N_1028[0] ;
    output n11079;
    input n5712;
    input n5711;
    input n5710;
    input VCC_net;
    output n5212;
    output n5525;
    input n5817;
    input n5618;
    input n5617;
    output tx_uart_active_flag;
    output n4715;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n5591, n3, n1, n3982;
    wire [2:0]r_Bit_Index_c;   // src/uart_tx.v(33[16:27])
    wire [2:0]n312;
    
    wire n8063, n3_adj_1363;
    wire [9:0]n45;
    wire [9:0]r_Clock_Count;   // src/uart_tx.v(32[16:29])
    
    wire n10349, n10348, n10347, n10346, n10345, n10344, n10343, 
        n10342, n10341, n4, n8, n7, n3981, n11586, n11646, o_Tx_Serial_N_1057, 
        n11643, n11583;
    
    SB_LUT4 i9988_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_1025[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n5591));
    defparam i9988_4_lut.LUT_INIT = 16'h4445;
    SB_DFFE o_Tx_Serial_44 (.Q(UART_TX_c), .C(SLM_CLK_c), .E(n1), .D(n3));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(SLM_CLK_c), .D(n3982), 
            .R(r_SM_Main[2]));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(SLM_CLK_c), .D(n11691));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i1539_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index_c[1]), 
            .I2(r_Bit_Index_c[2]), .I3(GND_net), .O(n312[2]));
    defparam i1539_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index_c[1]), 
            .I2(r_Bit_Index_c[2]), .I3(GND_net), .O(n8063));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(SLM_CLK_c), .D(n5716));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(SLM_CLK_c), .D(n5715));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(SLM_CLK_c), .D(n5714));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(SLM_CLK_c), .D(n5713));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i9920_4_lut_4_lut (.I0(\r_SM_Main_2__N_1025[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_1028[0] ), .O(n11079));   // src/uart_tx.v(41[7] 140[14])
    defparam i9920_4_lut_4_lut.LUT_INIT = 16'h8380;
    SB_DFF r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(SLM_CLK_c), .D(n5712));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i2908_2_lut_3_lut (.I0(\r_SM_Main_2__N_1025[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_1363));   // src/uart_tx.v(41[7] 140[14])
    defparam i2908_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 r_Clock_Count_1351_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[9]), .I3(n10349), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1351_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1351_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n10348), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1351_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(SLM_CLK_c), .D(n5711));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(SLM_CLK_c), .D(n5710));   // src/uart_tx.v(38[10] 141[8])
    SB_CARRY r_Clock_Count_1351_add_4_10 (.CI(n10348), .I0(GND_net), .I1(r_Clock_Count[8]), 
            .CO(n10349));
    SB_LUT4 r_Clock_Count_1351_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n10347), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1351_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1351_add_4_9 (.CI(n10347), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n10348));
    SB_LUT4 r_Clock_Count_1351_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n10346), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1351_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1351_add_4_8 (.CI(n10346), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n10347));
    SB_LUT4 r_Clock_Count_1351_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n10345), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1351_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1351_add_4_7 (.CI(n10345), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n10346));
    SB_LUT4 r_Clock_Count_1351_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n10344), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1351_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1351_add_4_6 (.CI(n10344), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n10345));
    SB_LUT4 r_Clock_Count_1351_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n10343), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1351_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1351_add_4_5 (.CI(n10343), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n10344));
    SB_LUT4 r_Clock_Count_1351_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n10342), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1351_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1351_add_4_4 (.CI(n10342), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n10343));
    SB_LUT4 r_Clock_Count_1351_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n10341), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1351_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1351_add_4_3 (.CI(n10341), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n10342));
    SB_LUT4 r_Clock_Count_1351_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
<<<<<<< HEAD
    defparam r_Clock_Count_1351_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(SLM_CLK_c), .D(n3_adj_1363), 
            .R(r_SM_Main[2]));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index_c[1]), .C(SLM_CLK_c), .E(n5212), 
            .D(n312[1]), .R(n5525));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index_c[2]), .C(SLM_CLK_c), .E(n5212), 
            .D(n312[2]), .R(n5525));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i4066_3_lut (.I0(n5212), .I1(n8063), .I2(r_SM_Main[1]), .I3(GND_net), 
            .O(n5525));   // src/uart_tx.v(38[10] 141[8])
    defparam i4066_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1532_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n312[1]));   // src/uart_tx.v(96[36:51])
    defparam i1532_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY r_Clock_Count_1351_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n10341));
=======
    defparam r_Clock_Count_1193_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n10214));
    SB_DFFESR r_Clock_Count_1193__i9 (.Q(r_Clock_Count[9]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[9]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i8 (.Q(r_Clock_Count[8]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[8]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i7 (.Q(r_Clock_Count[7]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[7]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i6 (.Q(r_Clock_Count[6]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[6]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i5 (.Q(r_Clock_Count[5]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[5]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i4 (.Q(r_Clock_Count[4]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[4]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i3 (.Q(r_Clock_Count[3]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[3]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i2 (.Q(r_Clock_Count[2]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[2]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i1 (.Q(r_Clock_Count[1]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[1]), .R(n4797));   // src/uart_tx.v(116[34:51])
    SB_LUT4 i10362_4_lut_4_lut (.I0(\r_SM_Main_2__N_841[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_844[0] ), .O(n10805));
    defparam i10362_4_lut_4_lut.LUT_INIT = 16'h8380;
    SB_LUT4 i2385_2_lut_3_lut (.I0(\r_SM_Main_2__N_841[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_1));
    defparam i2385_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_DFF r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(SLM_CLK_c), .D(n4890));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Active_46 (.Q(tx_uart_active_flag), .C(SLM_CLK_c), .D(n4889));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(SLM_CLK_c), .D(n5192));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(SLM_CLK_c), .D(n5191));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(SLM_CLK_c), .D(n5190));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(SLM_CLK_c), .D(n5189));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(SLM_CLK_c), .D(n5187));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i10392_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_841[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n4797));
    defparam i10392_4_lut.LUT_INIT = 16'h4445;
    SB_DFF r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(SLM_CLK_c), .D(n5171));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(SLM_CLK_c), .D(n5170));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(SLM_CLK_c), .E(n10955), 
            .D(n312[1]), .R(n10961));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(SLM_CLK_c), .E(n10955), 
            .D(n312[2]), .R(n10961));   // src/uart_tx.v(38[10] 141[8])
=======
module \uart_tx(CLKS_PER_BIT=20)  (GND_net, VCC_net, UART_TX_c, SLM_CLK_c, 
            r_SM_Main, \r_SM_Main_2__N_1026[1] , \r_Bit_Index[0] , n6966, 
            r_Tx_Data, n6965, n6964, n6963, n6962, n6961, n6960, 
            n6950, n16231, n5024, n5460, \r_SM_Main_2__N_1029[0] , 
            n4314, n5576, n5575, tx_uart_active_flag, n4) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    output UART_TX_c;
    input SLM_CLK_c;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_1026[1] ;
    output \r_Bit_Index[0] ;
    input n6966;
    output [7:0]r_Tx_Data;
    input n6965;
    input n6964;
    input n6963;
    input n6962;
    input n6961;
    input n6960;
    input n6950;
    input n16231;
    output n5024;
    output n5460;
    input \r_SM_Main_2__N_1029[0] ;
    output n4314;
    input n5576;
    input n5575;
    output tx_uart_active_flag;
    output n4;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [9:0]n45;
    wire [9:0]r_Clock_Count;   // src/uart_tx.v(32[16:29])
    
    wire n3, n1, n3602, n12196, n5541;
    wire [2:0]r_Bit_Index;   // src/uart_tx.v(33[16:27])
    wire [2:0]n312;
    
    wire n9003, n3_adj_1363, n4_c, n8, n7, n3601, n15160, n15136, 
        o_Tx_Serial_N_1058, n15157, n15133, n12204, n12203, n12202, 
        n12201, n12200, n12199, n12198, n12197;
    
    SB_LUT4 r_Clock_Count_1441_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1441_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFE o_Tx_Serial_44 (.Q(UART_TX_c), .C(SLM_CLK_c), .E(n1), .D(n3));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(SLM_CLK_c), .D(n3602), 
            .R(r_SM_Main[2]));   // src/uart_tx.v(38[10] 141[8])
    SB_CARRY r_Clock_Count_1441_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n12196));
    SB_LUT4 i12348_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_1026[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n5541));
    defparam i12348_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1622_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n312[1]));   // src/uart_tx.v(96[36:51])
    defparam i1622_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(SLM_CLK_c), .D(n6966));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(SLM_CLK_c), .D(n6965));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(SLM_CLK_c), .D(n6964));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(SLM_CLK_c), .D(n6963));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(SLM_CLK_c), .D(n6962));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(SLM_CLK_c), .D(n6961));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(SLM_CLK_c), .D(n6960));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFE r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n6950));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(SLM_CLK_c), .D(n16231));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i1629_2_lut_3_lut (.I0(\r_Bit_Index[0] ), .I1(r_Bit_Index[1]), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n312[2]));
    defparam i1629_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(SLM_CLK_c), .E(n5024), 
            .D(n312[2]), .R(n5460));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(SLM_CLK_c), .E(n5024), 
            .D(n312[1]), .R(n5460));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i2_2_lut_3_lut (.I0(\r_Bit_Index[0] ), .I1(r_Bit_Index[1]), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n9003));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFFESR r_Clock_Count_1441__i0 (.Q(r_Clock_Count[0]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[0]), .R(n5541));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1441__i9 (.Q(r_Clock_Count[9]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[9]), .R(n5541));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1441__i8 (.Q(r_Clock_Count[8]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[8]), .R(n5541));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1441__i7 (.Q(r_Clock_Count[7]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[7]), .R(n5541));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1441__i6 (.Q(r_Clock_Count[6]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[6]), .R(n5541));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1441__i5 (.Q(r_Clock_Count[5]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[5]), .R(n5541));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1441__i4 (.Q(r_Clock_Count[4]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[4]), .R(n5541));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1441__i3 (.Q(r_Clock_Count[3]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[3]), .R(n5541));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1441__i2 (.Q(r_Clock_Count[2]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[2]), .R(n5541));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1441__i1 (.Q(r_Clock_Count[1]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[1]), .R(n5541));   // src/uart_tx.v(116[34:51])
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_1026[1] ), .O(n5024));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_1029[0] ), .O(n4314));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(SLM_CLK_c), .D(n3_adj_1363), 
            .R(r_SM_Main[2]));   // src/uart_tx.v(38[10] 141[8])
>>>>>>> Stashed changes
>>>>>>> master
    SB_LUT4 i1_3_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[1]), 
            .I3(GND_net), .O(n4_c));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i2_2_lut (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[9]), .I2(GND_net), 
            .I3(GND_net), .O(n8));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[6]), .I2(r_Clock_Count[4]), 
            .I3(n4_c), .O(n7));
    defparam i1_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i5_4_lut (.I0(r_Clock_Count[5]), .I1(n7), .I2(r_Clock_Count[8]), 
<<<<<<< HEAD
            .I3(n8), .O(\r_SM_Main_2__N_1025[1] ));
=======
<<<<<<< Updated upstream
            .I3(n8), .O(\r_SM_Main_2__N_841[1] ));
>>>>>>> master
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2531_4_lut (.I0(\r_SM_Main_2__N_1028[0] ), .I1(n8063), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_1025[1] ), .O(n3981));   // src/uart_tx.v(41[7] 140[14])
    defparam i2531_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i2532_3_lut (.I0(n3981), .I1(\r_SM_Main_2__N_1025[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n3982));   // src/uart_tx.v(41[7] 140[14])
    defparam i2532_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i670925_i1_3_lut (.I0(n11586), .I1(n11646), .I2(r_Bit_Index_c[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_1057));
    defparam i670925_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_55_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_1057), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // src/uart_tx.v(41[7] 140[14])
    defparam r_SM_Main_2__I_0_55_i3_3_lut.LUT_INIT = 16'he5e5;
<<<<<<< HEAD
    SB_DFFESR r_Clock_Count_1351__i1 (.Q(r_Clock_Count[1]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[1]), .R(n5591));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1351__i2 (.Q(r_Clock_Count[2]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[2]), .R(n5591));   // src/uart_tx.v(116[34:51])
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_1025[1] ), .O(n5212));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_DFFESR r_Clock_Count_1351__i3 (.Q(r_Clock_Count[3]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[3]), .R(n5591));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1351__i4 (.Q(r_Clock_Count[4]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[4]), .R(n5591));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1351__i5 (.Q(r_Clock_Count[5]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[5]), .R(n5591));   // src/uart_tx.v(116[34:51])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n5817));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(SLM_CLK_c), .D(n5618));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Active_46 (.Q(tx_uart_active_flag), .C(SLM_CLK_c), .D(n5617));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_1028[0] ), .O(n4715));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index_c[1]), .O(n11643));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFFESR r_Clock_Count_1351__i6 (.Q(r_Clock_Count[6]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[6]), .R(n5591));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1351__i7 (.Q(r_Clock_Count[7]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[7]), .R(n5591));   // src/uart_tx.v(116[34:51])
    SB_LUT4 n11643_bdd_4_lut (.I0(n11643), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index_c[1]), .O(n11646));
    defparam n11643_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR r_Clock_Count_1351__i8 (.Q(r_Clock_Count[8]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[8]), .R(n5591));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1351__i9 (.Q(r_Clock_Count[9]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[9]), .R(n5591));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1351__i0 (.Q(r_Clock_Count[0]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[0]), .R(n5591));   // src/uart_tx.v(116[34:51])
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_10052 (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index_c[1]), .O(n11583));
    defparam r_Bit_Index_0__bdd_4_lut_10052.LUT_INIT = 16'he4aa;
    SB_LUT4 n11583_bdd_4_lut (.I0(n11583), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index_c[1]), .O(n11586));
    defparam n11583_bdd_4_lut.LUT_INIT = 16'haad8;
=======
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(n7576));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n11099), 
            .I2(n11100), .I3(r_Bit_Index[2]), .O(n12803));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n12803_bdd_4_lut (.I0(n12803), .I1(n11082), .I2(n11081), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_873));
    defparam n12803_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1365_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n312[1]));   // src/uart_tx.v(96[36:51])
    defparam i1365_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9261_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n11099));
    defparam i9261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9262_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n11100));
    defparam i9262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9244_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n11082));
    defparam i9244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9243_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n11081));
    defparam i9243_3_lut.LUT_INIT = 16'hcaca;
=======
            .I3(n8), .O(\r_SM_Main_2__N_1026[1] ));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2142_4_lut (.I0(\r_SM_Main_2__N_1029[0] ), .I1(n9003), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_1026[1] ), .O(n3601));   // src/uart_tx.v(41[7] 140[14])
    defparam i2142_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i2143_3_lut (.I0(n3601), .I1(\r_SM_Main_2__N_1026[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n3602));   // src/uart_tx.v(41[7] 140[14])
    defparam i2143_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7997244_i1_3_lut (.I0(n15160), .I1(n15136), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_1058));
    defparam i7997244_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_55_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_1058), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // src/uart_tx.v(41[7] 140[14])
    defparam r_SM_Main_2__I_0_55_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n15157));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n15157_bdd_4_lut (.I0(n15157), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n15160));
    defparam n15157_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_12931 (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n15133));
    defparam r_Bit_Index_0__bdd_4_lut_12931.LUT_INIT = 16'he4aa;
    SB_LUT4 n15133_bdd_4_lut (.I0(n15133), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n15136));
    defparam n15133_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(SLM_CLK_c), .D(n5576));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Active_46 (.Q(tx_uart_active_flag), .C(SLM_CLK_c), .D(n5575));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i12284_4_lut_4_lut (.I0(\r_SM_Main_2__N_1026[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_1029[0] ), .O(n4));   // src/uart_tx.v(41[7] 140[14])
    defparam i12284_4_lut_4_lut.LUT_INIT = 16'h8380;
    SB_LUT4 i2781_2_lut_3_lut (.I0(\r_SM_Main_2__N_1026[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_1363));   // src/uart_tx.v(41[7] 140[14])
    defparam i2781_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 r_Clock_Count_1441_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[9]), .I3(n12204), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1441_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1441_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n12203), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1441_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1441_add_4_10 (.CI(n12203), .I0(GND_net), .I1(r_Clock_Count[8]), 
            .CO(n12204));
    SB_LUT4 r_Clock_Count_1441_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n12202), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1441_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1441_add_4_9 (.CI(n12202), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n12203));
    SB_LUT4 r_Clock_Count_1441_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n12201), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1441_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1441_add_4_8 (.CI(n12201), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n12202));
    SB_LUT4 r_Clock_Count_1441_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n12200), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1441_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1441_add_4_7 (.CI(n12200), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n12201));
    SB_LUT4 r_Clock_Count_1441_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n12199), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1441_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1441_add_4_6 (.CI(n12199), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n12200));
    SB_LUT4 i3986_3_lut (.I0(n5024), .I1(n9003), .I2(r_SM_Main[1]), .I3(GND_net), 
            .O(n5460));   // src/uart_tx.v(38[10] 141[8])
    defparam i3986_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 r_Clock_Count_1441_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n12198), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1441_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1441_add_4_5 (.CI(n12198), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n12199));
    SB_LUT4 r_Clock_Count_1441_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n12197), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1441_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1441_add_4_4 (.CI(n12197), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n12198));
    SB_LUT4 r_Clock_Count_1441_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n12196), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1441_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1441_add_4_3 (.CI(n12196), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n12197));
>>>>>>> Stashed changes
>>>>>>> master
    
endmodule
//
// Verilog Description of module fifo_dc_32_lut_gen2
//

<<<<<<< HEAD
module fifo_dc_32_lut_gen2 (n30, n31, n5731, \REG.mem_28_0 , FIFO_CLK_c, 
            GND_net, n5726, \REG.mem_27_0 , n5725, \REG.mem_26_0 , 
            rd_fifo_en_w, DEBUG_5_c_0, SLM_CLK_c, DEBUG_1_c, reset_per_frame, 
            n5723, \REG.mem_25_0 , \REG.mem_16_0 , \REG.mem_17_0 , \rd_addr_r[0] , 
            \REG.mem_18_0 , \REG.mem_19_0 , n5721, \REG.mem_24_0 , \rd_grey_sync_r[0] , 
            \wr_addr_r[4] , DEBUG_9_c, wr_grey_sync_r, n5719, \REG.mem_23_0 , 
            \aempty_flag_impl.ae_flag_nxt_w , DEBUG_6_c, VCC_net, n5718, 
            \REG.mem_22_0 , n5717, \REG.mem_21_0 , dc32_fifo_full, \REG.mem_20_0 , 
            \rd_addr_nxt_c_5__N_572[2] , n5708, n5707, \REG.mem_14_0 , 
            \REG.mem_15_0 , \REG.mem_13_0 , \REG.mem_12_0 , n5691, rp_sync1_r, 
            n5690, n5689, n5688, n5687, n5686, n5685, n5684, n5683, 
            n5682, n5681, n5679, n7, n6, \REG.mem_2_0 , \REG.mem_3_0 , 
            \REG.mem_1_0 , \REG.mem_0_0 , n5677, \rd_addr_r[5] , n5675, 
            wp_sync1_r, n5674, n5673, n5672, n5671, \rd_grey_sync_r[4] , 
            \rd_grey_sync_r[3] , \rd_grey_sync_r[2] , \rd_grey_sync_r[1] , 
            n5670, n5669, n5668, n5667, n5666, n59, n47, n5664, 
            n5663, n5662, n5661, \wr_addr_nxt_c[0] , \wr_addr_nxt_c[1] , 
            n5659, \rd_addr_p1_w[0] , n5657, n5655, \REG.mem_6_0 , 
            \REG.mem_7_0 , dc32_fifo_read_enable, n5645, \REG.mem_11_0 , 
            \REG.mem_30_0 , \REG.mem_31_0 , \REG.mem_29_0 , \REG.mem_5_0 , 
            \REG.mem_4_0 , n5642, \REG.mem_10_0 , n5641, \REG.mem_9_0 , 
            n5640, \REG.mem_8_0 , \wr_addr_nxt_c[2] , \wr_addr_nxt_c[3] , 
            \wr_addr_nxt_c[4] , n25, \wr_grey_w[5] , n5639, dc32_fifo_write_enable, 
            n5638, n5637, n5635, n5634, n26, n5631, n5626, n5625, 
            n5624, n5623, n5622, n5615, n5611, \rd_addr_nxt_c_5__N_572[4] , 
            n5766, n5607, n24, n5762, n22, n20, n5751, n5750, 
            n5749, n23, n21, n5742, n28, n34, n35, n5735, n32, 
            n33, n29, n27) /* synthesis syn_module_defined=1 */ ;
    output n30;
    output n31;
    input n5731;
    output \REG.mem_28_0 ;
=======
<<<<<<< Updated upstream
module usb3_if (reset_per_frame, reset_per_frame_latched, SLM_CLK_c, DEBUG_3_c, 
            DEBUG_2_c, FIFO_CLK_c, \dc32_fifo_data_in[0] , DEBUG_5_c, 
            buffer_switch_done, buffer_switch_done_latched, VCC_net, FT_OE_c, 
            n571, GND_net, n575, write_to_dc32_fifo_latched_N_425, n2352, 
            n4911, n4910, n4907, FIFO_D15_c_15, FIFO_D14_c_14, FIFO_D13_c_13, 
            FIFO_D12_c_12, FIFO_D11_c_11, FIFO_D10_c_10, FIFO_D9_c_9, 
            FIFO_D8_c_8, FIFO_D7_c_7, FIFO_D6_c_6, FIFO_D5_c_5, FIFO_D4_c_4, 
            FIFO_D3_c_3, FIFO_D2_c_2, FIFO_D1_c_1, dc32_fifo_almost_full, 
            \dc32_fifo_data_in[15] , \dc32_fifo_data_in[14] , \dc32_fifo_data_in[13] , 
            \dc32_fifo_data_in[12] , \dc32_fifo_data_in[11] , \dc32_fifo_data_in[10] , 
            \dc32_fifo_data_in[9] , \dc32_fifo_data_in[8] , \dc32_fifo_data_in[7] , 
            \dc32_fifo_data_in[6] , \dc32_fifo_data_in[5] , \dc32_fifo_data_in[4] , 
            \dc32_fifo_data_in[3] , \dc32_fifo_data_in[2] , \dc32_fifo_data_in[1] , 
            DEBUG_1_c_c, FT_OE_N_420) /* synthesis syn_module_defined=1 */ ;
    input reset_per_frame;
    output reset_per_frame_latched;
    input SLM_CLK_c;
    input DEBUG_3_c;
    output DEBUG_2_c;
>>>>>>> master
    input FIFO_CLK_c;
    input GND_net;
    input n5726;
    output \REG.mem_27_0 ;
    input n5725;
    output \REG.mem_26_0 ;
    output rd_fifo_en_w;
    output DEBUG_5_c_0;
    input SLM_CLK_c;
    output DEBUG_1_c;
    input reset_per_frame;
    input n5723;
    output \REG.mem_25_0 ;
    output \REG.mem_16_0 ;
    output \REG.mem_17_0 ;
    output \rd_addr_r[0] ;
    output \REG.mem_18_0 ;
    output \REG.mem_19_0 ;
    input n5721;
    output \REG.mem_24_0 ;
    output \rd_grey_sync_r[0] ;
    output \wr_addr_r[4] ;
    output DEBUG_9_c;
    output [5:0]wr_grey_sync_r;
    input n5719;
    output \REG.mem_23_0 ;
    input \aempty_flag_impl.ae_flag_nxt_w ;
    output DEBUG_6_c;
    input VCC_net;
    input n5718;
    output \REG.mem_22_0 ;
    input n5717;
    output \REG.mem_21_0 ;
    output dc32_fifo_full;
    output \REG.mem_20_0 ;
    output \rd_addr_nxt_c_5__N_572[2] ;
    input n5708;
    input n5707;
    output \REG.mem_14_0 ;
    output \REG.mem_15_0 ;
    output \REG.mem_13_0 ;
    output \REG.mem_12_0 ;
    input n5691;
    output [5:0]rp_sync1_r;
    input n5690;
    input n5689;
    input n5688;
    input n5687;
    input n5686;
    input n5685;
    input n5684;
    input n5683;
    input n5682;
    input n5681;
    input n5679;
    output n7;
    output n6;
    output \REG.mem_2_0 ;
    output \REG.mem_3_0 ;
    output \REG.mem_1_0 ;
    output \REG.mem_0_0 ;
    input n5677;
    output \rd_addr_r[5] ;
    input n5675;
    output [5:0]wp_sync1_r;
    input n5674;
    input n5673;
    input n5672;
    input n5671;
    output \rd_grey_sync_r[4] ;
    output \rd_grey_sync_r[3] ;
    output \rd_grey_sync_r[2] ;
    output \rd_grey_sync_r[1] ;
    input n5670;
    input n5669;
    input n5668;
    input n5667;
    input n5666;
    output n59;
    input n47;
    input n5664;
    input n5663;
    input n5662;
    input n5661;
    output \wr_addr_nxt_c[0] ;
    output \wr_addr_nxt_c[1] ;
    input n5659;
    output \rd_addr_p1_w[0] ;
    input n5657;
    input n5655;
    output \REG.mem_6_0 ;
    output \REG.mem_7_0 ;
    input dc32_fifo_read_enable;
    input n5645;
    output \REG.mem_11_0 ;
    output \REG.mem_30_0 ;
    output \REG.mem_31_0 ;
    output \REG.mem_29_0 ;
    output \REG.mem_5_0 ;
    output \REG.mem_4_0 ;
    input n5642;
    output \REG.mem_10_0 ;
    input n5641;
    output \REG.mem_9_0 ;
    input n5640;
    output \REG.mem_8_0 ;
    output \wr_addr_nxt_c[2] ;
    output \wr_addr_nxt_c[3] ;
    output \wr_addr_nxt_c[4] ;
    output n25;
    output \wr_grey_w[5] ;
    input n5639;
    input dc32_fifo_write_enable;
    input n5638;
    input n5637;
    input n5635;
    input n5634;
    output n26;
    input n5631;
    input n5626;
    input n5625;
    input n5624;
    input n5623;
    input n5622;
    input n5615;
    input n5611;
    output \rd_addr_nxt_c_5__N_572[4] ;
    input n5766;
    input n5607;
    output n24;
    input n5762;
    output n22;
    output n20;
    input n5751;
    input n5750;
    input n5749;
    output n23;
    output n21;
    input n5742;
    output n28;
    output n34;
    output n35;
    input n5735;
    output n32;
    output n33;
    output n29;
    output n27;
    
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1 lscc_fifo_dc_inst (.n30(n30), 
            .n31(n31), .n5731(n5731), .\REG.mem_28_0 (\REG.mem_28_0 ), 
            .FIFO_CLK_c(FIFO_CLK_c), .GND_net(GND_net), .n5726(n5726), 
            .\REG.mem_27_0 (\REG.mem_27_0 ), .n5725(n5725), .\REG.mem_26_0 (\REG.mem_26_0 ), 
            .rd_fifo_en_w(rd_fifo_en_w), .DEBUG_5_c_0(DEBUG_5_c_0), .SLM_CLK_c(SLM_CLK_c), 
            .DEBUG_1_c(DEBUG_1_c), .reset_per_frame(reset_per_frame), .n5723(n5723), 
            .\REG.mem_25_0 (\REG.mem_25_0 ), .\REG.mem_16_0 (\REG.mem_16_0 ), 
            .\REG.mem_17_0 (\REG.mem_17_0 ), .rd_addr_r({Open_2, Open_3, 
            Open_4, Open_5, Open_6, \rd_addr_r[0] }), .\REG.mem_18_0 (\REG.mem_18_0 ), 
            .\REG.mem_19_0 (\REG.mem_19_0 ), .n5721(n5721), .\REG.mem_24_0 (\REG.mem_24_0 ), 
            .\rd_grey_sync_r[0] (\rd_grey_sync_r[0] ), .\wr_addr_r[4] (\wr_addr_r[4] ), 
            .DEBUG_9_c(DEBUG_9_c), .wr_grey_sync_r({wr_grey_sync_r}), .n5719(n5719), 
            .\REG.mem_23_0 (\REG.mem_23_0 ), .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .DEBUG_6_c(DEBUG_6_c), .VCC_net(VCC_net), .n5718(n5718), .\REG.mem_22_0 (\REG.mem_22_0 ), 
            .n5717(n5717), .\REG.mem_21_0 (\REG.mem_21_0 ), .dc32_fifo_full(dc32_fifo_full), 
            .\REG.mem_20_0 (\REG.mem_20_0 ), .\rd_addr_nxt_c_5__N_572[2] (\rd_addr_nxt_c_5__N_572[2] ), 
            .n5708(n5708), .n5707(n5707), .\REG.mem_14_0 (\REG.mem_14_0 ), 
            .\REG.mem_15_0 (\REG.mem_15_0 ), .\REG.mem_13_0 (\REG.mem_13_0 ), 
            .\REG.mem_12_0 (\REG.mem_12_0 ), .n5691(n5691), .rp_sync1_r({rp_sync1_r}), 
            .n5690(n5690), .n5689(n5689), .n5688(n5688), .n5687(n5687), 
            .n5686(n5686), .n5685(n5685), .n5684(n5684), .n5683(n5683), 
            .n5682(n5682), .n5681(n5681), .n5679(n5679), .n7(n7), .n6(n6), 
            .\REG.mem_2_0 (\REG.mem_2_0 ), .\REG.mem_3_0 (\REG.mem_3_0 ), 
            .\REG.mem_1_0 (\REG.mem_1_0 ), .\REG.mem_0_0 (\REG.mem_0_0 ), 
            .n5677(n5677), .\rd_addr_r[5] (\rd_addr_r[5] ), .n5675(n5675), 
            .wp_sync1_r({wp_sync1_r}), .n5674(n5674), .n5673(n5673), .n5672(n5672), 
            .n5671(n5671), .\rd_grey_sync_r[4] (\rd_grey_sync_r[4] ), .\rd_grey_sync_r[3] (\rd_grey_sync_r[3] ), 
            .\rd_grey_sync_r[2] (\rd_grey_sync_r[2] ), .\rd_grey_sync_r[1] (\rd_grey_sync_r[1] ), 
            .n5670(n5670), .n5669(n5669), .n5668(n5668), .n5667(n5667), 
            .n5666(n5666), .n59(n59), .n47(n47), .n5664(n5664), .n5663(n5663), 
            .n5662(n5662), .n5661(n5661), .\wr_addr_nxt_c[0] (\wr_addr_nxt_c[0] ), 
            .\wr_addr_nxt_c[1] (\wr_addr_nxt_c[1] ), .n5659(n5659), .\rd_addr_p1_w[0] (\rd_addr_p1_w[0] ), 
            .n5657(n5657), .n5655(n5655), .\REG.mem_6_0 (\REG.mem_6_0 ), 
            .\REG.mem_7_0 (\REG.mem_7_0 ), .dc32_fifo_read_enable(dc32_fifo_read_enable), 
            .n5645(n5645), .\REG.mem_11_0 (\REG.mem_11_0 ), .\REG.mem_30_0 (\REG.mem_30_0 ), 
            .\REG.mem_31_0 (\REG.mem_31_0 ), .\REG.mem_29_0 (\REG.mem_29_0 ), 
            .\REG.mem_5_0 (\REG.mem_5_0 ), .\REG.mem_4_0 (\REG.mem_4_0 ), 
            .n5642(n5642), .\REG.mem_10_0 (\REG.mem_10_0 ), .n5641(n5641), 
            .\REG.mem_9_0 (\REG.mem_9_0 ), .n5640(n5640), .\REG.mem_8_0 (\REG.mem_8_0 ), 
            .\wr_addr_nxt_c[2] (\wr_addr_nxt_c[2] ), .\wr_addr_nxt_c[3] (\wr_addr_nxt_c[3] ), 
            .\wr_addr_nxt_c[4] (\wr_addr_nxt_c[4] ), .n25(n25), .\wr_grey_w[5] (\wr_grey_w[5] ), 
            .n5639(n5639), .dc32_fifo_write_enable(dc32_fifo_write_enable), 
            .n5638(n5638), .n5637(n5637), .n5635(n5635), .n5634(n5634), 
            .n26(n26), .n5631(n5631), .n5626(n5626), .n5625(n5625), 
            .n5624(n5624), .n5623(n5623), .n5622(n5622), .n5615(n5615), 
            .n5611(n5611), .\rd_addr_nxt_c_5__N_572[4] (\rd_addr_nxt_c_5__N_572[4] ), 
            .n5766(n5766), .n5607(n5607), .n24(n24), .n5762(n5762), 
            .n22(n22), .n20(n20), .n5751(n5751), .n5750(n5750), .n5749(n5749), 
            .n23(n23), .n21(n21), .n5742(n5742), .n28(n28), .n34(n34), 
            .n35(n35), .n5735(n5735), .n32(n32), .n33(n33), .n29(n29), 
            .n27(n27)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_dc_32_lut_gen.v(53[33] 72[34])
    
endmodule
//
// Verilog Description of module fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1
//

module fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1 (n30, 
            n31, n5731, \REG.mem_28_0 , FIFO_CLK_c, GND_net, n5726, 
            \REG.mem_27_0 , n5725, \REG.mem_26_0 , rd_fifo_en_w, DEBUG_5_c_0, 
            SLM_CLK_c, DEBUG_1_c, reset_per_frame, n5723, \REG.mem_25_0 , 
            \REG.mem_16_0 , \REG.mem_17_0 , rd_addr_r, \REG.mem_18_0 , 
            \REG.mem_19_0 , n5721, \REG.mem_24_0 , \rd_grey_sync_r[0] , 
            \wr_addr_r[4] , DEBUG_9_c, wr_grey_sync_r, n5719, \REG.mem_23_0 , 
            \aempty_flag_impl.ae_flag_nxt_w , DEBUG_6_c, VCC_net, n5718, 
            \REG.mem_22_0 , n5717, \REG.mem_21_0 , dc32_fifo_full, \REG.mem_20_0 , 
            \rd_addr_nxt_c_5__N_572[2] , n5708, n5707, \REG.mem_14_0 , 
            \REG.mem_15_0 , \REG.mem_13_0 , \REG.mem_12_0 , n5691, rp_sync1_r, 
            n5690, n5689, n5688, n5687, n5686, n5685, n5684, n5683, 
            n5682, n5681, n5679, n7, n6, \REG.mem_2_0 , \REG.mem_3_0 , 
            \REG.mem_1_0 , \REG.mem_0_0 , n5677, \rd_addr_r[5] , n5675, 
            wp_sync1_r, n5674, n5673, n5672, n5671, \rd_grey_sync_r[4] , 
            \rd_grey_sync_r[3] , \rd_grey_sync_r[2] , \rd_grey_sync_r[1] , 
            n5670, n5669, n5668, n5667, n5666, n59, n47, n5664, 
            n5663, n5662, n5661, \wr_addr_nxt_c[0] , \wr_addr_nxt_c[1] , 
            n5659, \rd_addr_p1_w[0] , n5657, n5655, \REG.mem_6_0 , 
            \REG.mem_7_0 , dc32_fifo_read_enable, n5645, \REG.mem_11_0 , 
            \REG.mem_30_0 , \REG.mem_31_0 , \REG.mem_29_0 , \REG.mem_5_0 , 
            \REG.mem_4_0 , n5642, \REG.mem_10_0 , n5641, \REG.mem_9_0 , 
            n5640, \REG.mem_8_0 , \wr_addr_nxt_c[2] , \wr_addr_nxt_c[3] , 
            \wr_addr_nxt_c[4] , n25, \wr_grey_w[5] , n5639, dc32_fifo_write_enable, 
            n5638, n5637, n5635, n5634, n26, n5631, n5626, n5625, 
            n5624, n5623, n5622, n5615, n5611, \rd_addr_nxt_c_5__N_572[4] , 
            n5766, n5607, n24, n5762, n22, n20, n5751, n5750, 
            n5749, n23, n21, n5742, n28, n34, n35, n5735, n32, 
            n33, n29, n27) /* synthesis syn_module_defined=1 */ ;
    output n30;
    output n31;
    input n5731;
    output \REG.mem_28_0 ;
    input FIFO_CLK_c;
    input GND_net;
    input n5726;
    output \REG.mem_27_0 ;
    input n5725;
    output \REG.mem_26_0 ;
    output rd_fifo_en_w;
    output DEBUG_5_c_0;
    input SLM_CLK_c;
    output DEBUG_1_c;
    input reset_per_frame;
    input n5723;
    output \REG.mem_25_0 ;
    output \REG.mem_16_0 ;
    output \REG.mem_17_0 ;
    output [5:0]rd_addr_r;
    output \REG.mem_18_0 ;
    output \REG.mem_19_0 ;
    input n5721;
    output \REG.mem_24_0 ;
    output \rd_grey_sync_r[0] ;
    output \wr_addr_r[4] ;
    output DEBUG_9_c;
    output [5:0]wr_grey_sync_r;
    input n5719;
    output \REG.mem_23_0 ;
    input \aempty_flag_impl.ae_flag_nxt_w ;
    output DEBUG_6_c;
    input VCC_net;
    input n5718;
    output \REG.mem_22_0 ;
    input n5717;
    output \REG.mem_21_0 ;
    output dc32_fifo_full;
    output \REG.mem_20_0 ;
    output \rd_addr_nxt_c_5__N_572[2] ;
    input n5708;
    input n5707;
    output \REG.mem_14_0 ;
    output \REG.mem_15_0 ;
    output \REG.mem_13_0 ;
    output \REG.mem_12_0 ;
    input n5691;
    output [5:0]rp_sync1_r;
    input n5690;
    input n5689;
    input n5688;
    input n5687;
    input n5686;
    input n5685;
    input n5684;
    input n5683;
    input n5682;
    input n5681;
    input n5679;
    output n7;
    output n6;
    output \REG.mem_2_0 ;
    output \REG.mem_3_0 ;
    output \REG.mem_1_0 ;
    output \REG.mem_0_0 ;
    input n5677;
    output \rd_addr_r[5] ;
    input n5675;
    output [5:0]wp_sync1_r;
    input n5674;
    input n5673;
    input n5672;
    input n5671;
    output \rd_grey_sync_r[4] ;
    output \rd_grey_sync_r[3] ;
    output \rd_grey_sync_r[2] ;
    output \rd_grey_sync_r[1] ;
    input n5670;
    input n5669;
    input n5668;
    input n5667;
    input n5666;
    output n59;
    input n47;
    input n5664;
    input n5663;
    input n5662;
    input n5661;
    output \wr_addr_nxt_c[0] ;
    output \wr_addr_nxt_c[1] ;
    input n5659;
    output \rd_addr_p1_w[0] ;
    input n5657;
    input n5655;
    output \REG.mem_6_0 ;
    output \REG.mem_7_0 ;
    input dc32_fifo_read_enable;
    input n5645;
    output \REG.mem_11_0 ;
    output \REG.mem_30_0 ;
    output \REG.mem_31_0 ;
    output \REG.mem_29_0 ;
    output \REG.mem_5_0 ;
    output \REG.mem_4_0 ;
    input n5642;
    output \REG.mem_10_0 ;
    input n5641;
    output \REG.mem_9_0 ;
    input n5640;
    output \REG.mem_8_0 ;
    output \wr_addr_nxt_c[2] ;
    output \wr_addr_nxt_c[3] ;
    output \wr_addr_nxt_c[4] ;
    output n25;
    output \wr_grey_w[5] ;
    input n5639;
    input dc32_fifo_write_enable;
    input n5638;
    input n5637;
    input n5635;
    input n5634;
    output n26;
    input n5631;
    input n5626;
    input n5625;
    input n5624;
    input n5623;
    input n5622;
    input n5615;
    input n5611;
    output \rd_addr_nxt_c_5__N_572[4] ;
    input n5766;
    input n5607;
    output n24;
    input n5762;
    output n22;
    output n20;
    input n5751;
    input n5750;
    input n5749;
    output n23;
    output n21;
    input n5742;
    output n28;
    output n34;
    output n35;
    input n5735;
    output n32;
    output n33;
    output n29;
    output n27;
    
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n6_c;
    wire [5:0]wr_addr_r;   // src/fifo_dc_32_lut_gen.v(196[29:38])
    
    wire n10298, n10299;
    wire [31:0]rd_data_o_31__N_597;
    
    wire \afull_flag_impl.af_flag_nxt_w ;
    wire [5:0]wr_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(200[30:42])
    
    wire n10297, n11329, n11330, n10296;
    wire [5:0]rp_sync2_r;   // src/fifo_dc_32_lut_gen.v(202[37:47])
    wire [5:0]rp_sync_w;   // src/fifo_dc_32_lut_gen.v(205[30:39])
    wire [5:0]rd_grey_w;   // src/fifo_dc_32_lut_gen.v(224[38:47])
    
    wire n8, n11157, n11211, n11169, empty_nxt_c_N_635, n11221;
    wire [5:0]wr_grey_w;   // src/fifo_dc_32_lut_gen.v(203[38:47])
    
    wire n11350, n11267, n11619, n11598, n11604;
    wire [5:0]rd_addr_r_c;   // src/fifo_dc_32_lut_gen.v(217[29:38])
    
    wire n11622, full_nxt_c_N_632, n11336, n11335;
    wire [5:0]rd_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(221[30:42])
    
    wire n5680;
    wire [5:0]rd_addr_nxt_c_5__N_572;
    
    wire n11685, n11328;
    wire [5:0]wp_sync2_r;   // src/fifo_dc_32_lut_gen.v(223[37:47])
    wire [5:0]n1;
    
    wire n10249;
    wire [5:0]rd_sig_diff0_w;   // src/fifo_dc_32_lut_gen.v(233[30:44])
    wire [5:0]wp_sync_w;   // src/fifo_dc_32_lut_gen.v(226[30:39])
    
    wire n10248, n11601, n5678, n10247, n5676, n10246;
    wire [5:0]n1_adj_1362;
    
    wire n10285, n10375, n8_adj_1354, n10284, n6_adj_1355, n10245, 
        n73, n7_adj_1358, n10283;
    wire [5:0]wr_sig_diff0_w;   // src/fifo_dc_32_lut_gen.v(212[30:44])
    
    wire n5047, n11183, n11217, n8_adj_1359, n7_adj_1360, n11595, 
        n9, n11265, n10418, n11667, n11670, n10282, n11649, n10281, 
        n8069, n7_adj_1361, n11652, n11634, n11333, n10305, n11334, 
        n10304, n10303, n10302, n10301, n11589, n11592, n10300, 
        n11631;
    
    SB_LUT4 EnabledDecoder_2_i30_2_lut_3_lut_4_lut (.I0(n6_c), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[2]), .O(n30));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i30_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i31_2_lut_3_lut_4_lut (.I0(n6_c), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[2]), .O(n31));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i31_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_DFF i2726_2727 (.Q(\REG.mem_28_0 ), .C(FIFO_CLK_c), .D(n5731));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY wr_addr_r_5__I_0_128_5 (.CI(n10298), .I0(wr_addr_r[3]), .I1(GND_net), 
            .CO(n10299));
    SB_DFF i2630_2631 (.Q(\REG.mem_27_0 ), .C(FIFO_CLK_c), .D(n5726));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2534_2535 (.Q(\REG.mem_26_0 ), .C(FIFO_CLK_c), .D(n5725));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFE \REG.out_raw__i1  (.Q(DEBUG_5_c_0), .C(SLM_CLK_c), .E(rd_fifo_en_w), 
            .D(rd_data_o_31__N_597[0]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFSR \afull_flag_impl.af_flag_ext_r_111  (.Q(DEBUG_1_c), .C(FIFO_CLK_c), 
            .D(\afull_flag_impl.af_flag_nxt_w ), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(410[29] 422[32])
    SB_LUT4 wr_addr_r_5__I_0_128_4_lut (.I0(GND_net), .I1(wr_addr_r[2]), 
            .I2(GND_net), .I3(n10297), .O(wr_addr_p1_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF i2438_2439 (.Q(\REG.mem_25_0 ), .C(FIFO_CLK_c), .D(n5723));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY wr_addr_r_5__I_0_128_4 (.CI(n10297), .I0(wr_addr_r[2]), .I1(GND_net), 
            .CO(n10298));
    SB_LUT4 i9749_3_lut (.I0(\REG.mem_16_0 ), .I1(\REG.mem_17_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11329));
    defparam i9749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9750_3_lut (.I0(\REG.mem_18_0 ), .I1(\REG.mem_19_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11330));
    defparam i9750_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2342_2343 (.Q(\REG.mem_24_0 ), .C(FIFO_CLK_c), .D(n5721));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wr_addr_r_5__I_0_128_3_lut (.I0(GND_net), .I1(wr_addr_r[1]), 
            .I2(GND_net), .I3(n10296), .O(wr_addr_p1_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rp_sync2_r_5__I_0_124_i1_2_lut (.I0(rp_sync2_r[4]), .I1(rp_sync2_r[5]), 
            .I2(GND_net), .I3(GND_net), .O(rp_sync_w[4]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam rp_sync2_r_5__I_0_124_i1_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut (.I0(rp_sync2_r[0]), .I1(rp_sync_w[1]), .I2(GND_net), 
            .I3(GND_net), .O(rp_sync_w[0]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
<<<<<<< HEAD
    SB_LUT4 i2_3_lut (.I0(rp_sync2_r[3]), .I1(rp_sync2_r[4]), .I2(rp_sync2_r[5]), 
            .I3(GND_net), .O(rp_sync_w[3]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i2_3_lut.LUT_INIT = 16'h6969;
    SB_CARRY wr_addr_r_5__I_0_128_3 (.CI(n10296), .I0(wr_addr_r[1]), .I1(GND_net), 
            .CO(n10297));
    SB_LUT4 i1_2_lut_adj_36 (.I0(rp_sync2_r[2]), .I1(rp_sync_w[3]), .I2(GND_net), 
            .I3(GND_net), .O(rp_sync_w[2]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_adj_36.LUT_INIT = 16'h6666;
    SB_DFFSR rd_grey_sync_r__i0 (.Q(\rd_grey_sync_r[0] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[0]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_LUT4 i2_4_lut (.I0(wr_addr_p1_w[2]), .I1(wr_addr_p1_w[5]), .I2(rp_sync_w[2]), 
            .I3(rp_sync2_r[5]), .O(n8));
    defparam i2_4_lut.LUT_INIT = 16'h1248;
    SB_LUT4 i9581_4_lut (.I0(wr_addr_p1_w[3]), .I1(wr_addr_p1_w[0]), .I2(rp_sync_w[3]), 
            .I3(rp_sync_w[0]), .O(n11157));
    defparam i9581_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 i9634_4_lut (.I0(wr_addr_p1_w[4]), .I1(wr_addr_p1_w[1]), .I2(rp_sync_w[4]), 
            .I3(rp_sync_w[1]), .O(n11211));
    defparam i9634_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 i9593_4_lut (.I0(wr_addr_r[1]), .I1(\wr_addr_r[4] ), .I2(rp_sync_w[1]), 
            .I3(rp_sync_w[4]), .O(n11169));
    defparam i9593_4_lut.LUT_INIT = 16'hedb7;
    SB_DFFSS empty_ext_r_114 (.Q(DEBUG_9_c), .C(SLM_CLK_c), .D(empty_nxt_c_N_635), 
            .S(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_LUT4 i9644_4_lut (.I0(wr_addr_r[3]), .I1(wr_addr_r[0]), .I2(rp_sync_w[3]), 
            .I3(rp_sync_w[0]), .O(n11221));
    defparam i9644_4_lut.LUT_INIT = 16'hedb7;
    SB_DFFSR wr_grey_sync_r__i0 (.Q(wr_grey_sync_r[0]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[0]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_LUT4 i9859_3_lut (.I0(n11211), .I1(n11157), .I2(n8), .I3(GND_net), 
            .O(n11350));   // src/fifo_dc_32_lut_gen.v(300[45:114])
    defparam i9859_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i9689_4_lut (.I0(n11221), .I1(wr_addr_r[2]), .I2(n11169), 
            .I3(rp_sync_w[2]), .O(n11267));
    defparam i9689_4_lut.LUT_INIT = 16'hfefb;
    SB_DFF i2246_2247 (.Q(\REG.mem_23_0 ), .C(FIFO_CLK_c), .D(n5719));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFS \aempty_flag_impl.ae_flag_ext_r_120  (.Q(DEBUG_6_c), .C(SLM_CLK_c), 
            .D(\aempty_flag_impl.ae_flag_nxt_w ), .S(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(669[37] 672[40])
    SB_LUT4 wr_addr_r_5__I_0_128_2_lut (.I0(GND_net), .I1(wr_addr_r[0]), 
            .I2(GND_net), .I3(VCC_net), .O(wr_addr_p1_w[0])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF i2150_2151 (.Q(\REG.mem_22_0 ), .C(FIFO_CLK_c), .D(n5718));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2054_2055 (.Q(\REG.mem_21_0 ), .C(FIFO_CLK_c), .D(n5717));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY wr_addr_r_5__I_0_128_2 (.CI(VCC_net), .I0(wr_addr_r[0]), .I1(GND_net), 
            .CO(n10296));
    SB_LUT4 n11619_bdd_4_lut (.I0(n11619), .I1(n11598), .I2(n11604), .I3(rd_addr_r_c[3]), 
            .O(n11622));
    defparam n11619_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR full_ext_r_107 (.Q(dc32_fifo_full), .C(FIFO_CLK_c), .D(full_nxt_c_N_632), 
            .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 i9756_3_lut (.I0(\REG.mem_22_0 ), .I1(\REG.mem_23_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11336));
    defparam i9756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9755_3_lut (.I0(\REG.mem_20_0 ), .I1(\REG.mem_21_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11335));
    defparam i9755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_nxt_c_5__I_0_138_i2_2_lut_4_lut (.I0(rd_addr_r_c[1]), 
            .I1(rd_addr_p1_w[1]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_5__N_572[2] ), 
            .O(rd_grey_w[1]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_5__I_0_138_i2_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4221_2_lut_4_lut (.I0(rd_addr_r_c[1]), .I1(rd_addr_p1_w[1]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n5680));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4221_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 rd_addr_nxt_c_5__I_0_138_i1_2_lut_4_lut (.I0(rd_addr_r_c[1]), 
            .I1(rd_addr_p1_w[1]), .I2(rd_fifo_en_w), .I3(rd_addr_nxt_c_5__N_572[0]), 
            .O(rd_grey_w[0]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_5__I_0_138_i1_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_DFF i1958_1959 (.Q(\REG.mem_20_0 ), .C(FIFO_CLK_c), .D(n5708));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1862_1863 (.Q(\REG.mem_19_0 ), .C(FIFO_CLK_c), .D(n5707));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut (.I0(rd_addr_r[0]), .I1(\REG.mem_14_0 ), 
            .I2(\REG.mem_15_0 ), .I3(rd_addr_r_c[1]), .O(n11685));
    defparam rd_addr_r_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n11685_bdd_4_lut (.I0(n11685), .I1(\REG.mem_13_0 ), .I2(\REG.mem_12_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11328));
    defparam n11685_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF rp_sync1_r__i1 (.Q(rp_sync1_r[1]), .C(FIFO_CLK_c), .D(n5691));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i2 (.Q(rp_sync1_r[2]), .C(FIFO_CLK_c), .D(n5690));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i3 (.Q(rp_sync1_r[3]), .C(FIFO_CLK_c), .D(n5689));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i4 (.Q(rp_sync1_r[4]), .C(FIFO_CLK_c), .D(n5688));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i5 (.Q(rp_sync1_r[5]), .C(FIFO_CLK_c), .D(n5687));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF i1766_1767 (.Q(\REG.mem_18_0 ), .C(FIFO_CLK_c), .D(n5686));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync2_r__i1 (.Q(rp_sync2_r[1]), .C(FIFO_CLK_c), .D(n5685));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i2 (.Q(rp_sync2_r[2]), .C(FIFO_CLK_c), .D(n5684));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i3 (.Q(rp_sync2_r[3]), .C(FIFO_CLK_c), .D(n5683));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i4 (.Q(rp_sync2_r[4]), .C(FIFO_CLK_c), .D(n5682));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i5 (.Q(rp_sync2_r[5]), .C(FIFO_CLK_c), .D(n5681));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rd_addr_r__i1 (.Q(rd_addr_r_c[1]), .C(SLM_CLK_c), .D(n5680));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i2 (.Q(rd_addr_r_c[2]), .C(SLM_CLK_c), .D(n5679));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_7_lut (.I0(rd_sig_diff0_w[2]), .I1(wp_sync2_r[5]), 
            .I2(n1[5]), .I3(n10249), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_7_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_6_lut (.I0(rd_sig_diff0_w[3]), .I1(wp_sync_w[4]), 
            .I2(n1[4]), .I3(n10248), .O(n6)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_6_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10042 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_0 ), 
            .I2(\REG.mem_3_0 ), .I3(rd_addr_r_c[1]), .O(n11601));
    defparam rd_addr_r_0__bdd_4_lut_10042.LUT_INIT = 16'he4aa;
    SB_DFF rd_addr_r__i3 (.Q(rd_addr_r_c[3]), .C(SLM_CLK_c), .D(n5678));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_LUT4 n11601_bdd_4_lut (.I0(n11601), .I1(\REG.mem_1_0 ), .I2(\REG.mem_0_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11604));
    defparam n11601_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY wp_sync2_r_5__I_0_135_add_2_6 (.CI(n10248), .I0(wp_sync_w[4]), 
            .I1(n1[4]), .CO(n10249));
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_5_lut (.I0(GND_net), .I1(wp_sync_w[3]), 
            .I2(n1[3]), .I3(n10247), .O(rd_sig_diff0_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF rd_addr_r__i4 (.Q(rd_addr_r_c[4]), .C(SLM_CLK_c), .D(n5677));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i5 (.Q(\rd_addr_r[5] ), .C(SLM_CLK_c), .D(n5676));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_CARRY wp_sync2_r_5__I_0_135_add_2_5 (.CI(n10247), .I0(wp_sync_w[3]), 
            .I1(n1[3]), .CO(n10248));
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_4_lut (.I0(GND_net), .I1(wp_sync_w[2]), 
            .I2(n1[2]), .I3(n10246), .O(rd_sig_diff0_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF wp_sync1_r__i1 (.Q(wp_sync1_r[1]), .C(SLM_CLK_c), .D(n5675));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_CARRY wp_sync2_r_5__I_0_135_add_2_4 (.CI(n10246), .I0(wp_sync_w[2]), 
            .I1(n1[2]), .CO(n10247));
    SB_LUT4 wr_addr_r_5__I_0_add_2_7_lut (.I0(n10375), .I1(wr_grey_sync_r[5]), 
            .I2(n1_adj_1362[5]), .I3(n10285), .O(\afull_flag_impl.af_flag_nxt_w )) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_7_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 wr_addr_r_5__I_0_add_2_6_lut (.I0(n6_adj_1355), .I1(\wr_addr_r[4] ), 
            .I2(rp_sync_w[4]), .I3(n10284), .O(n8_adj_1354)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_6_lut.LUT_INIT = 16'h8228;
    SB_DFFSR wr_grey_sync_r__i4 (.Q(wr_grey_sync_r[4]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[4]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFSR wr_grey_sync_r__i3 (.Q(wr_grey_sync_r[3]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[3]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFSR wr_grey_sync_r__i2 (.Q(wr_grey_sync_r[2]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[2]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFSR wr_grey_sync_r__i1 (.Q(wr_grey_sync_r[1]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[1]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFF wp_sync1_r__i2 (.Q(wp_sync1_r[2]), .C(SLM_CLK_c), .D(n5674));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i3 (.Q(wp_sync1_r[3]), .C(SLM_CLK_c), .D(n5673));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i4 (.Q(wp_sync1_r[4]), .C(SLM_CLK_c), .D(n5672));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i5 (.Q(wp_sync1_r[5]), .C(SLM_CLK_c), .D(n5671));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFFSR rd_grey_sync_r__i4 (.Q(\rd_grey_sync_r[4] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[4]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i3 (.Q(\rd_grey_sync_r[3] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[3]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i2 (.Q(\rd_grey_sync_r[2] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[2]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i1 (.Q(\rd_grey_sync_r[1] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[1]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFF wp_sync2_r__i1 (.Q(wp_sync2_r[1]), .C(SLM_CLK_c), .D(n5670));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i2 (.Q(wp_sync2_r[2]), .C(SLM_CLK_c), .D(n5669));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i3 (.Q(wp_sync2_r[3]), .C(SLM_CLK_c), .D(n5668));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i4 (.Q(wp_sync2_r[4]), .C(SLM_CLK_c), .D(n5667));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i5 (.Q(wp_sync2_r[5]), .C(SLM_CLK_c), .D(n5666));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_3_lut (.I0(n73), .I1(wp_sync_w[1]), 
            .I2(n1[1]), .I3(n10245), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY wp_sync2_r_5__I_0_135_add_2_3 (.CI(n10245), .I0(wp_sync_w[1]), 
            .I1(n1[1]), .CO(n10246));
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_2_lut (.I0(n47), .I1(wp_sync_w[0]), 
            .I2(n1[0]), .I3(VCC_net), .O(n73)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY wp_sync2_r_5__I_0_135_add_2_2 (.CI(VCC_net), .I0(wp_sync_w[0]), 
            .I1(n1[0]), .CO(n10245));
    SB_DFF i1670_1671 (.Q(\REG.mem_17_0 ), .C(FIFO_CLK_c), .D(n5664));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wr_grey_sync_r__i5 (.Q(wr_grey_sync_r[5]), .C(FIFO_CLK_c), .D(n5663));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_CARRY wr_addr_r_5__I_0_add_2_6 (.CI(n10284), .I0(\wr_addr_r[4] ), 
            .I1(rp_sync_w[4]), .CO(n10285));
    SB_LUT4 wr_addr_r_5__I_0_add_2_5_lut (.I0(wr_sig_diff0_w[2]), .I1(wr_addr_r[3]), 
            .I2(rp_sync_w[3]), .I3(n10283), .O(n7_adj_1358)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_5_lut.LUT_INIT = 16'h8228;
    SB_DFF i1574_1575 (.Q(\REG.mem_16_0 ), .C(FIFO_CLK_c), .D(n5662));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1478_1479 (.Q(\REG.mem_15_0 ), .C(FIFO_CLK_c), .D(n5661));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wr_addr_nxt_c_5__I_0_136_i1_2_lut (.I0(\wr_addr_nxt_c[0] ), .I1(\wr_addr_nxt_c[1] ), 
            .I2(GND_net), .I3(GND_net), .O(wr_grey_w[0]));   // src/fifo_dc_32_lut_gen.v(253[28:66])
    defparam wr_addr_nxt_c_5__I_0_136_i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_37 (.I0(wp_sync2_r[5]), .I1(wp_sync2_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5047));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_37.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_38 (.I0(wp_sync2_r[1]), .I1(wp_sync_w[2]), .I2(GND_net), 
            .I3(GND_net), .O(wp_sync_w[1]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_38.LUT_INIT = 16'h6666;
    SB_LUT4 i9607_4_lut (.I0(rd_addr_r_c[3]), .I1(rd_addr_r[0]), .I2(wp_sync_w[3]), 
            .I3(wp_sync_w[0]), .O(n11183));
    defparam i9607_4_lut.LUT_INIT = 16'h7bde;
    SB_DFF i1382_1383 (.Q(\REG.mem_14_0 ), .C(FIFO_CLK_c), .D(n5659));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9640_4_lut (.I0(rd_addr_r_c[2]), .I1(rd_addr_r_c[4]), .I2(wp_sync_w[2]), 
            .I3(n5047), .O(n11217));
    defparam i9640_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut_adj_39 (.I0(wp_sync2_r[5]), .I1(rd_addr_p1_w[1]), .I2(rd_addr_p1_w[5]), 
            .I3(wp_sync_w[1]), .O(n8_adj_1359));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i2_4_lut_adj_39.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut (.I0(rd_addr_p1_w[2]), .I1(\rd_addr_p1_w[0] ), .I2(wp_sync_w[2]), 
            .I3(wp_sync_w[0]), .O(n7_adj_1360));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i1_4_lut.LUT_INIT = 16'h7bde;
    SB_DFF i1286_1287 (.Q(\REG.mem_13_0 ), .C(FIFO_CLK_c), .D(n5657));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1190_1191 (.Q(\REG.mem_12_0 ), .C(FIFO_CLK_c), .D(n5655));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10019 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_0 ), 
            .I2(\REG.mem_7_0 ), .I3(rd_addr_r_c[1]), .O(n11595));
    defparam rd_addr_r_0__bdd_4_lut_10019.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut (.I0(rd_addr_p1_w[3]), .I1(rd_addr_p1_w[4]), .I2(wp_sync_w[3]), 
            .I3(n5047), .O(n9));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i3_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i9687_4_lut (.I0(n11217), .I1(rd_addr_r_c[1]), .I2(n11183), 
            .I3(wp_sync_w[1]), .O(n11265));
    defparam i9687_4_lut.LUT_INIT = 16'hfbfe;
    SB_LUT4 i5_3_lut (.I0(n9), .I1(n7_adj_1360), .I2(n8_adj_1359), .I3(GND_net), 
            .O(n10418));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 empty_nxt_c_I_11_4_lut (.I0(n10418), .I1(n11265), .I2(DEBUG_9_c), 
            .I3(dc32_fifo_read_enable), .O(empty_nxt_c_N_635));   // src/fifo_dc_32_lut_gen.v(555[46:103])
    defparam empty_nxt_c_I_11_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 rd_addr_r_5__I_0_i1_3_lut (.I0(rd_addr_r[0]), .I1(\rd_addr_p1_w[0] ), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(rd_addr_nxt_c_5__N_572[0]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_5__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i1_1_lut (.I0(rd_addr_r[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_DFF i1094_1095 (.Q(\REG.mem_11_0 ), .C(FIFO_CLK_c), .D(n5645));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10086 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_0 ), 
            .I2(\REG.mem_31_0 ), .I3(rd_addr_r_c[1]), .O(n11667));
    defparam rd_addr_r_0__bdd_4_lut_10086.LUT_INIT = 16'he4aa;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i2_1_lut (.I0(rd_addr_r_c[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n11667_bdd_4_lut (.I0(n11667), .I1(\REG.mem_29_0 ), .I2(\REG.mem_28_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11670));
    defparam n11667_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY wr_addr_r_5__I_0_add_2_5 (.CI(n10283), .I0(wr_addr_r[3]), .I1(rp_sync_w[3]), 
            .CO(n10284));
    SB_LUT4 wr_addr_r_5__I_0_add_2_4_lut (.I0(GND_net), .I1(wr_addr_r[2]), 
            .I2(rp_sync_w[2]), .I3(n10282), .O(wr_sig_diff0_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11595_bdd_4_lut (.I0(n11595), .I1(\REG.mem_5_0 ), .I2(\REG.mem_4_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11598));
    defparam n11595_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i998_999 (.Q(\REG.mem_10_0 ), .C(FIFO_CLK_c), .D(n5642));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i902_903 (.Q(\REG.mem_9_0 ), .C(FIFO_CLK_c), .D(n5641));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i806_807 (.Q(\REG.mem_8_0 ), .C(FIFO_CLK_c), .D(n5640));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut (.I0(rd_addr_r_c[1]), .I1(n11335), .I2(n11336), 
            .I3(rd_addr_r_c[2]), .O(n11649));
    defparam rd_addr_r_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_CARRY wr_addr_r_5__I_0_add_2_4 (.CI(n10282), .I0(wr_addr_r[2]), .I1(rp_sync_w[2]), 
            .CO(n10283));
    SB_LUT4 wr_addr_r_5__I_0_add_2_3_lut (.I0(n8069), .I1(wr_addr_r[1]), 
            .I2(rp_sync_w[1]), .I3(n10281), .O(n6_adj_1355)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY wr_addr_r_5__I_0_add_2_3 (.CI(n10281), .I0(wr_addr_r[1]), .I1(rp_sync_w[1]), 
            .CO(n10282));
    SB_LUT4 wr_addr_nxt_c_5__I_0_136_i2_2_lut (.I0(\wr_addr_nxt_c[1] ), .I1(\wr_addr_nxt_c[2] ), 
            .I2(GND_net), .I3(GND_net), .O(wr_grey_w[1]));   // src/fifo_dc_32_lut_gen.v(253[28:66])
    defparam wr_addr_nxt_c_5__I_0_136_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 wr_addr_nxt_c_5__I_0_136_i3_2_lut (.I0(\wr_addr_nxt_c[2] ), .I1(\wr_addr_nxt_c[3] ), 
            .I2(GND_net), .I3(GND_net), .O(wr_grey_w[2]));   // src/fifo_dc_32_lut_gen.v(253[28:66])
    defparam wr_addr_nxt_c_5__I_0_136_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 wr_addr_nxt_c_5__I_0_136_i4_2_lut (.I0(\wr_addr_nxt_c[3] ), .I1(\wr_addr_nxt_c[4] ), 
            .I2(GND_net), .I3(GND_net), .O(wr_grey_w[3]));   // src/fifo_dc_32_lut_gen.v(253[28:66])
    defparam wr_addr_nxt_c_5__I_0_136_i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 EnabledDecoder_2_i25_2_lut_4_lut (.I0(n7_adj_1361), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[3]), .O(n25));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i25_2_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 wr_addr_nxt_c_5__I_0_136_i5_2_lut (.I0(\wr_addr_nxt_c[4] ), .I1(\wr_grey_w[5] ), 
            .I2(GND_net), .I3(GND_net), .O(wr_grey_w[4]));   // src/fifo_dc_32_lut_gen.v(253[28:66])
    defparam wr_addr_nxt_c_5__I_0_136_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n11649_bdd_4_lut (.I0(n11649), .I1(n11330), .I2(n11329), .I3(rd_addr_r_c[2]), 
            .O(n11652));
    defparam n11649_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(wp_sync2_r[2]), .I1(wp_sync2_r[3]), 
            .I2(wp_sync2_r[5]), .I3(wp_sync2_r[4]), .O(wp_sync_w[2]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut (.I0(n7_adj_1358), .I1(n8_adj_1354), .I2(GND_net), 
            .I3(GND_net), .O(n10375));
    defparam i4_2_lut.LUT_INIT = 16'h8888;
    SB_DFF i710_711 (.Q(\REG.mem_7_0 ), .C(FIFO_CLK_c), .D(n5639));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wr_addr_r_5__I_0_inv_0_i6_1_lut (.I0(rp_sync2_r[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1362[5]));   // src/fifo_dc_32_lut_gen.v(212[47:78])
    defparam wr_addr_r_5__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 wr_addr_r_5__I_0_add_2_2_lut (.I0(dc32_fifo_write_enable), .I1(wr_addr_r[0]), 
            .I2(rp_sync_w[0]), .I3(VCC_net), .O(n8069)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_DFF i614_615 (.Q(\REG.mem_6_0 ), .C(FIFO_CLK_c), .D(n5638));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY wr_addr_r_5__I_0_add_2_2 (.CI(VCC_net), .I0(wr_addr_r[0]), 
            .I1(rp_sync_w[0]), .CO(n10281));
    SB_DFF i518_519 (.Q(\REG.mem_5_0 ), .C(FIFO_CLK_c), .D(n5637));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_en_i_I_0_2_lut (.I0(dc32_fifo_read_enable), .I1(DEBUG_9_c), 
            .I2(GND_net), .I3(GND_net), .O(rd_fifo_en_w));   // src/fifo_dc_32_lut_gen.v(241[29:51])
    defparam rd_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_DFF i422_423 (.Q(\REG.mem_4_0 ), .C(FIFO_CLK_c), .D(n5635));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9753_3_lut (.I0(n11634), .I1(n11670), .I2(rd_addr_r_c[2]), 
            .I3(GND_net), .O(n11333));
    defparam i9753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_5__I_0_137_7_lut (.I0(GND_net), .I1(\rd_addr_r[5] ), 
            .I2(GND_net), .I3(n10305), .O(rd_addr_p1_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF i326_327 (.Q(\REG.mem_3_0 ), .C(FIFO_CLK_c), .D(n5634));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9754_3_lut (.I0(n11652), .I1(n11333), .I2(rd_addr_r_c[3]), 
            .I3(GND_net), .O(n11334));
    defparam i9754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_5__I_0_137_6_lut (.I0(GND_net), .I1(rd_addr_r_c[4]), 
            .I2(GND_net), .I3(n10304), .O(rd_addr_p1_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i670322_i1_3_lut (.I0(n11622), .I1(n11334), .I2(rd_addr_r_c[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_597[0]));
    defparam i670322_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i26_2_lut_4_lut (.I0(n6_c), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[3]), .O(n26));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i26_2_lut_4_lut.LUT_INIT = 16'h0800;
    SB_DFF i134_135 (.Q(\REG.mem_1_0 ), .C(FIFO_CLK_c), .D(n5631));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY rd_addr_r_5__I_0_137_6 (.CI(n10304), .I0(rd_addr_r_c[4]), .I1(GND_net), 
            .CO(n10305));
    SB_LUT4 rd_addr_r_5__I_0_137_5_lut (.I0(GND_net), .I1(rd_addr_r_c[3]), 
            .I2(GND_net), .I3(n10303), .O(rd_addr_p1_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rd_addr_r_5__I_0_137_5 (.CI(n10303), .I0(rd_addr_r_c[3]), .I1(GND_net), 
            .CO(n10304));
    SB_LUT4 rd_addr_r_5__I_0_137_4_lut (.I0(GND_net), .I1(rd_addr_r_c[2]), 
            .I2(GND_net), .I3(n10302), .O(rd_addr_p1_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rd_addr_r_5__I_0_137_4 (.CI(n10302), .I0(rd_addr_r_c[2]), .I1(GND_net), 
            .CO(n10303));
    SB_DFF wp_sync2_r__i0 (.Q(wp_sync2_r[0]), .C(SLM_CLK_c), .D(n5626));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_LUT4 rd_addr_r_5__I_0_137_3_lut (.I0(GND_net), .I1(rd_addr_r_c[1]), 
            .I2(GND_net), .I3(n10301), .O(rd_addr_p1_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF wp_sync1_r__i0 (.Q(wp_sync1_r[0]), .C(SLM_CLK_c), .D(n5625));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10014 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_0 ), 
            .I2(\REG.mem_11_0 ), .I3(rd_addr_r_c[1]), .O(n11589));
    defparam rd_addr_r_0__bdd_4_lut_10014.LUT_INIT = 16'he4aa;
    SB_DFF rd_addr_r__i0 (.Q(rd_addr_r[0]), .C(SLM_CLK_c), .D(n5624));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_LUT4 n11589_bdd_4_lut (.I0(n11589), .I1(\REG.mem_9_0 ), .I2(\REG.mem_8_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11592));
    defparam n11589_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY rd_addr_r_5__I_0_137_3 (.CI(n10301), .I0(rd_addr_r_c[1]), .I1(GND_net), 
            .CO(n10302));
    SB_DFF rp_sync2_r__i0 (.Q(rp_sync2_r[0]), .C(FIFO_CLK_c), .D(n5623));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_LUT4 rd_addr_r_5__I_0_137_2_lut (.I0(GND_net), .I1(rd_addr_r[0]), 
            .I2(GND_net), .I3(VCC_net), .O(\rd_addr_p1_w[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i3_1_lut (.I0(rd_addr_r_c[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_DFF rp_sync1_r__i0 (.Q(rp_sync1_r[0]), .C(FIFO_CLK_c), .D(n5622));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF i230_231 (.Q(\REG.mem_2_0 ), .C(FIFO_CLK_c), .D(n5615));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i38_39 (.Q(\REG.mem_0_0 ), .C(FIFO_CLK_c), .D(n5611));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_5__I_0_i5_3_lut (.I0(rd_addr_r_c[4]), .I1(rd_addr_p1_w[4]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_5__N_572[4] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_5__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i4_1_lut (.I0(rd_addr_r_c[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i5_1_lut (.I0(rd_addr_r_c[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 wp_sync2_r_5__I_0_130_i1_2_lut (.I0(wp_sync2_r[4]), .I1(wp_sync2_r[5]), 
            .I2(GND_net), .I3(GND_net), .O(wp_sync_w[4]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam wp_sync2_r_5__I_0_130_i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i6_1_lut (.I0(\rd_addr_r[5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rd_addr_r_5__I_0_i3_3_lut (.I0(rd_addr_r_c[2]), .I1(rd_addr_p1_w[2]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_5__N_572[2] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_5__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_5__I_0_123_i3_3_lut_4_lut (.I0(dc32_fifo_write_enable), 
            .I1(dc32_fifo_full), .I2(wr_addr_p1_w[2]), .I3(wr_addr_r[2]), 
            .O(\wr_addr_nxt_c[2] ));   // src/fifo_dc_32_lut_gen.v(240[29:50])
    defparam wr_addr_r_5__I_0_123_i3_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_addr_r_5__I_0_123_i4_3_lut_4_lut (.I0(dc32_fifo_write_enable), 
            .I1(dc32_fifo_full), .I2(wr_addr_p1_w[3]), .I3(wr_addr_r[3]), 
            .O(\wr_addr_nxt_c[3] ));   // src/fifo_dc_32_lut_gen.v(240[29:50])
    defparam wr_addr_r_5__I_0_123_i4_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3014_3015 (.Q(\REG.mem_31_0 ), .C(FIFO_CLK_c), .D(n5766));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wr_addr_r_5__I_0_123_i6_3_lut_4_lut (.I0(dc32_fifo_write_enable), 
            .I1(dc32_fifo_full), .I2(wr_addr_p1_w[5]), .I3(wr_grey_sync_r[5]), 
            .O(\wr_grey_w[5] ));   // src/fifo_dc_32_lut_gen.v(240[29:50])
    defparam wr_addr_r_5__I_0_123_i6_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF wr_addr_r__i0 (.Q(wr_addr_r[0]), .C(FIFO_CLK_c), .D(n5607));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 EnabledDecoder_2_i24_2_lut_4_lut (.I0(n7_adj_1361), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[3]), .O(n24));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i24_2_lut_4_lut.LUT_INIT = 16'h0800;
    SB_DFF i2918_2919 (.Q(\REG.mem_30_0 ), .C(FIFO_CLK_c), .D(n5762));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY rd_addr_r_5__I_0_137_2 (.CI(VCC_net), .I0(rd_addr_r[0]), .I1(GND_net), 
            .CO(n10301));
    SB_LUT4 EnabledDecoder_2_i22_2_lut_4_lut (.I0(n6_c), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[3]), .O(n22));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i22_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 wr_addr_r_5__I_0_123_i5_3_lut_4_lut (.I0(dc32_fifo_write_enable), 
            .I1(dc32_fifo_full), .I2(wr_addr_p1_w[4]), .I3(\wr_addr_r[4] ), 
            .O(\wr_addr_nxt_c[4] ));   // src/fifo_dc_32_lut_gen.v(240[29:50])
    defparam wr_addr_r_5__I_0_123_i5_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i20_2_lut_4_lut (.I0(n7_adj_1361), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[3]), .O(n20));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i20_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 wr_addr_r_5__I_0_128_7_lut (.I0(GND_net), .I1(wr_grey_sync_r[5]), 
            .I2(GND_net), .I3(n10300), .O(wr_addr_p1_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF wr_addr_r__i1 (.Q(wr_addr_r[1]), .C(FIFO_CLK_c), .D(n5751));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i2 (.Q(wr_addr_r[2]), .C(FIFO_CLK_c), .D(n5750));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 wr_addr_r_5__I_0_123_i1_3_lut_4_lut (.I0(dc32_fifo_write_enable), 
            .I1(dc32_fifo_full), .I2(wr_addr_p1_w[0]), .I3(wr_addr_r[0]), 
            .O(\wr_addr_nxt_c[0] ));   // src/fifo_dc_32_lut_gen.v(240[29:50])
    defparam wr_addr_r_5__I_0_123_i1_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF wr_addr_r__i3 (.Q(wr_addr_r[3]), .C(FIFO_CLK_c), .D(n5749));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 wr_addr_r_5__I_0_128_6_lut (.I0(GND_net), .I1(\wr_addr_r[4] ), 
            .I2(GND_net), .I3(n10299), .O(wr_addr_p1_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_5__I_0_128_6 (.CI(n10299), .I0(\wr_addr_r[4] ), .I1(GND_net), 
            .CO(n10300));
    SB_LUT4 EnabledDecoder_2_i23_2_lut_4_lut (.I0(n6_c), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[3]), .O(n23));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i23_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i21_2_lut_4_lut (.I0(n7_adj_1361), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[3]), .O(n21));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i21_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_DFF wr_addr_r__i4 (.Q(\wr_addr_r[4] ), .C(FIFO_CLK_c), .D(n5742));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 rd_addr_r_2__bdd_4_lut (.I0(rd_addr_r_c[2]), .I1(n11592), .I2(n11328), 
            .I3(rd_addr_r_c[3]), .O(n11619));
    defparam rd_addr_r_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i6_2_lut_3_lut (.I0(dc32_fifo_write_enable), 
            .I1(dc32_fifo_full), .I2(wr_addr_r[0]), .I3(GND_net), .O(n6_c));   // src/fifo_dc_32_lut_gen.v(240[29:50])
    defparam EnabledDecoder_2_i6_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1_2_lut_3_lut (.I0(wp_sync2_r[3]), .I1(wp_sync2_r[5]), .I2(wp_sync2_r[4]), 
            .I3(GND_net), .O(wp_sync_w[3]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 EnabledDecoder_2_i7_2_lut_3_lut (.I0(dc32_fifo_write_enable), 
            .I1(dc32_fifo_full), .I2(wr_addr_r[0]), .I3(GND_net), .O(n7_adj_1361));   // src/fifo_dc_32_lut_gen.v(240[29:50])
    defparam EnabledDecoder_2_i7_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_3_lut_adj_40 (.I0(wp_sync2_r[0]), .I1(wp_sync2_r[1]), 
            .I2(wp_sync_w[2]), .I3(GND_net), .O(wp_sync_w[0]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_adj_40.LUT_INIT = 16'h9696;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10071 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_0 ), 
            .I2(\REG.mem_27_0 ), .I3(rd_addr_r_c[1]), .O(n11631));
    defparam rd_addr_r_0__bdd_4_lut_10071.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i28_2_lut_4_lut (.I0(n7_adj_1361), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[3]), .O(n28));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i28_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i34_2_lut_3_lut_4_lut (.I0(n6_c), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[2]), .O(n34));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i34_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 EnabledDecoder_2_i35_2_lut_3_lut_4_lut (.I0(n6_c), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[2]), .O(n35));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i35_2_lut_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 wr_addr_r_5__I_0_123_i2_3_lut_4_lut (.I0(dc32_fifo_write_enable), 
            .I1(dc32_fifo_full), .I2(wr_addr_p1_w[1]), .I3(wr_addr_r[1]), 
            .O(\wr_addr_nxt_c[1] ));   // src/fifo_dc_32_lut_gen.v(240[29:50])
    defparam wr_addr_r_5__I_0_123_i2_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_nxt_c_5__I_0_138_i3_2_lut_4_lut (.I0(rd_addr_r_c[3]), 
            .I1(rd_addr_p1_w[3]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_5__N_572[2] ), 
            .O(rd_grey_w[2]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_5__I_0_138_i3_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 rd_addr_nxt_c_5__I_0_138_i4_2_lut_4_lut (.I0(rd_addr_r_c[3]), 
            .I1(rd_addr_p1_w[3]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_5__N_572[4] ), 
            .O(rd_grey_w[3]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_5__I_0_138_i4_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_DFF i2822_2823 (.Q(\REG.mem_29_0 ), .C(FIFO_CLK_c), .D(n5735));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n11631_bdd_4_lut (.I0(n11631), .I1(\REG.mem_25_0 ), .I2(\REG.mem_24_0 ), 
            .I3(rd_addr_r_c[1]), .O(n11634));
    defparam n11631_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4219_2_lut_4_lut (.I0(rd_addr_r_c[3]), .I1(rd_addr_p1_w[3]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n5678));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4219_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 wr_addr_r_5__I_0_128_5_lut (.I0(GND_net), .I1(wr_addr_r[3]), 
            .I2(GND_net), .I3(n10298), .O(wr_addr_p1_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_nxt_c_5__I_0_138_i5_2_lut_4_lut (.I0(\rd_addr_r[5] ), 
            .I1(rd_addr_p1_w[5]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_5__N_572[4] ), 
            .O(rd_grey_w[4]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_5__I_0_138_i5_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 full_nxt_c_I_10_4_lut_4_lut (.I0(dc32_fifo_write_enable), .I1(dc32_fifo_full), 
            .I2(n11350), .I3(n11267), .O(full_nxt_c_N_632));   // src/fifo_dc_32_lut_gen.v(240[29:50])
    defparam full_nxt_c_I_10_4_lut_4_lut.LUT_INIT = 16'h20ec;
    SB_LUT4 i4217_2_lut_4_lut (.I0(\rd_addr_r[5] ), .I1(rd_addr_p1_w[5]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n5676));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4217_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 EnabledDecoder_2_i32_2_lut_3_lut_4_lut (.I0(n7_adj_1361), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[2]), .O(n32));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i32_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 EnabledDecoder_2_i33_2_lut_3_lut_4_lut (.I0(n7_adj_1361), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[2]), .O(n33));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i33_2_lut_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i1_2_lut_3_lut_adj_41 (.I0(rp_sync2_r[2]), .I1(rp_sync_w[3]), 
            .I2(rp_sync2_r[1]), .I3(GND_net), .O(rp_sync_w[1]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_3_lut_adj_41.LUT_INIT = 16'h9696;
    SB_LUT4 EnabledDecoder_2_i29_2_lut_4_lut (.I0(n7_adj_1361), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[3]), .O(n29));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i29_2_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i27_2_lut_4_lut (.I0(n6_c), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[3]), .O(n27));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i27_2_lut_4_lut.LUT_INIT = 16'h0008;
=======
    SB_LUT4 i10447_3_lut (.I0(n10783), .I1(reset_per_frame_latched), .I2(n4181), 
            .I3(GND_net), .O(n4310));   // src/usb3_if.v(97[10] 190[8])
    defparam i10447_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_4_lut_adj_2 (.I0(n562[0]), .I1(n2266), .I2(n520), .I3(DEBUG_1_c_c), 
            .O(n10783));   // src/usb3_if.v(97[10] 190[8])
    defparam i1_4_lut_adj_2.LUT_INIT = 16'h0ace;
    SB_LUT4 i3306_4_lut (.I0(n4310), .I1(n562[2]), .I2(n562[0]), .I3(n2390), 
            .O(n4688));   // src/usb3_if.v(88[8] 191[4])
    defparam i3306_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 i1050_2_lut (.I0(n562[5]), .I1(dc32_fifo_almost_full), .I2(GND_net), 
            .I3(GND_net), .O(n2266));
    defparam i1050_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_1159_i3_4_lut (.I0(n2408), .I1(n3938), .I2(n2415), .I3(n1[0]), 
            .O(n2401));   // src/usb3_if.v(98[9] 189[16])
    defparam mux_1159_i3_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 mux_1159_i4_4_lut (.I0(n12077), .I1(n3942), .I2(n2415), .I3(n2408), 
            .O(n2402));   // src/usb3_if.v(98[9] 189[16])
    defparam mux_1159_i4_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i10300_2_lut (.I0(n21), .I1(dc32_fifo_empty_latched), .I2(GND_net), 
            .I3(GND_net), .O(n12077));   // src/usb3_if.v(98[9] 189[16])
    defparam i10300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i179_2_lut_3_lut (.I0(n524), .I1(dc32_fifo_almost_full), .I2(DEBUG_1_c_c), 
            .I3(GND_net), .O(n551));   // src/usb3_if.v(155[26] 157[24])
    defparam i179_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1647_3_lut_4_lut (.I0(n562[5]), .I1(n562[8]), .I2(n562[4]), 
            .I3(FT_OE_N_420), .O(n3014));   // src/usb3_if.v(98[9] 189[16])
    defparam i1647_3_lut_4_lut.LUT_INIT = 16'hfcfe;
    SB_LUT4 i10389_2_lut (.I0(n562[5]), .I1(reset_per_frame_latched), .I2(GND_net), 
            .I3(GND_net), .O(n2983));   // src/usb3_if.v(88[8] 191[4])
    defparam i10389_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_3_lut (.I0(n524), .I1(reset_per_frame_latched), .I2(n562[2]), 
            .I3(GND_net), .O(n4486));
    defparam i1_3_lut.LUT_INIT = 16'hdcdc;
    SB_LUT4 mux_1159_i1_4_lut (.I0(n12030), .I1(state_timeout_counter[0]), 
            .I2(n2415), .I3(n2408), .O(n2399));   // src/usb3_if.v(98[9] 189[16])
    defparam mux_1159_i1_4_lut.LUT_INIT = 16'h3a3f;
    SB_LUT4 i10282_2_lut (.I0(n21), .I1(dc32_fifo_empty_latched), .I2(GND_net), 
            .I3(GND_net), .O(n12030));   // src/usb3_if.v(98[9] 189[16])
    defparam i10282_2_lut.LUT_INIT = 16'h4444;
=======
module usb3_if (reset_per_frame, reset_per_frame_latched, SLM_CLK_c, dc32_fifo_empty, 
            VCC_net, FT_RD_c, FIFO_CLK_c, dc32_fifo_data_in, dc32_fifo_write_enable, 
            buffer_switch_done, buffer_switch_done_latched, GND_net, DEBUG_1_c, 
            n663, n7014, FR_RXF_c, FT_OE_c, DEBUG_3_c_0_c, FIFO_D1_c_1, 
            FIFO_D2_c_2, FIFO_D3_c_3, FIFO_D4_c_4, FIFO_D5_c_5, FIFO_D6_c_6, 
            FIFO_D7_c_7, FIFO_D8_c_8, FIFO_D9_c_9, FIFO_D10_c_10, FIFO_D11_c_11, 
            FIFO_D12_c_12, FIFO_D13_c_13, FIFO_D14_c_14, FIFO_D15_c_15, 
            FIFO_D16_c_16, FIFO_D17_c_17, FIFO_D18_c_18, FIFO_D19_c_19, 
            FIFO_D20_c_20, FIFO_D21_c_21, FIFO_D22_c_22, FIFO_D23_c_23, 
            FIFO_D24_c_24, FIFO_D25_c_25, FIFO_D26_c_26, FIFO_D27_c_27, 
            FIFO_D28_c_28, FIFO_D29_c_29, FIFO_D30_c_30, FIFO_D31_c_31) /* synthesis syn_module_defined=1 */ ;
    input reset_per_frame;
    output reset_per_frame_latched;
    input SLM_CLK_c;
    input dc32_fifo_empty;
    input VCC_net;
    output FT_RD_c;
    input FIFO_CLK_c;
    output [31:0]dc32_fifo_data_in;
    output dc32_fifo_write_enable;
    input buffer_switch_done;
    output buffer_switch_done_latched;
    input GND_net;
    input DEBUG_1_c;
    output n663;
    input n7014;
    input FR_RXF_c;
    output FT_OE_c;
    input DEBUG_3_c_0_c;
    input FIFO_D1_c_1;
    input FIFO_D2_c_2;
    input FIFO_D3_c_3;
    input FIFO_D4_c_4;
    input FIFO_D5_c_5;
    input FIFO_D6_c_6;
    input FIFO_D7_c_7;
    input FIFO_D8_c_8;
    input FIFO_D9_c_9;
    input FIFO_D10_c_10;
    input FIFO_D11_c_11;
    input FIFO_D12_c_12;
    input FIFO_D13_c_13;
    input FIFO_D14_c_14;
    input FIFO_D15_c_15;
    input FIFO_D16_c_16;
    input FIFO_D17_c_17;
    input FIFO_D18_c_18;
    input FIFO_D19_c_19;
    input FIFO_D20_c_20;
    input FIFO_D21_c_21;
    input FIFO_D22_c_22;
    input FIFO_D23_c_23;
    input FIFO_D24_c_24;
    input FIFO_D25_c_25;
    input FIFO_D26_c_26;
    input FIFO_D27_c_27;
    input FIFO_D28_c_28;
    input FIFO_D29_c_29;
    input FIFO_D30_c_30;
    input FIFO_D31_c_31;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    
    wire dc32_fifo_empty_latched, FT_RD_N_501;
    wire [31:0]dc32_fifo_data_in_latched;   // src/usb3_if.v(66[12:37])
    wire [15:0]n650;
    
    wire n4839, n5368, write_to_dc32_fifo_latched;
    wire [4:0]state_timeout_counter;   // src/usb3_if.v(64[11:32])
    
    wire n4454;
    wire [10:0]num_lines_clocked_out_10__N_441;
    wire [10:0]num_lines_clocked_out;   // src/usb3_if.v(63[12:33])
    
    wire n12115, n6, n12116, n3462;
    wire [31:0]n850;
    
    wire n5138, n5387, n12114, n2737, n2741, n8, n2727;
    wire [3:0]n187;
    
    wire n2744, n2726, n2725, n609, n4226, n605, FT_OE_N_491, 
        n12843, n10, n2724, write_to_dc32_fifo_latched_N_503, n3611;
    wire [6:0]n70;
    
    wire n5298;
    wire [5:0]num_words_curr_line_5__N_435;
    
    wire n4963, n5425, FT_OE_N_495, n172, n12877, n14301, n12113;
    wire [5:0]num_words_curr_line;   // src/usb3_if.v(60[11:30])
    
    wire n4772, n12112, n12111, n12110, n12109, n4983, n12108, 
        n8999, n11, n12107, n883, n18, n16, n20, n607, FT_OE_N_490, 
        n12121, n12120, n12119, n2723, n12840, n3458, n696, n3456, 
        n3452, n706, n709, n6_adj_1361, n6_adj_1362, n918, n8991, 
        n12118, n12117, n4757, n12270, n694, n3459, n8685;
    
    SB_DFF reset_per_frame_latched_109 (.Q(reset_per_frame_latched), .C(SLM_CLK_c), 
           .D(reset_per_frame));   // src/usb3_if.v(70[8] 83[4])
    SB_DFF dc32_fifo_empty_latched_110 (.Q(dc32_fifo_empty_latched), .C(SLM_CLK_c), 
           .D(dc32_fifo_empty));   // src/usb3_if.v(70[8] 83[4])
    SB_DFFESS FT_RD_112 (.Q(FT_RD_c), .C(FIFO_CLK_c), .E(VCC_net), .D(FT_RD_N_501), 
            .S(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFN dc32_fifo_data_in_i0 (.Q(dc32_fifo_data_in[0]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[0]));   // src/usb3_if.v(204[8] 207[4])
    SB_LUT4 i3894_4_lut_4_lut (.I0(n650[0]), .I1(n650[2]), .I2(n650[5]), 
            .I3(n4839), .O(n5368));
    defparam i3894_4_lut_4_lut.LUT_INIT = 16'h3200;
    SB_DFFN write_to_dc32_fifo_120 (.Q(dc32_fifo_write_enable), .C(FIFO_CLK_c), 
            .D(write_to_dc32_fifo_latched));   // src/usb3_if.v(204[8] 207[4])
    SB_DFF buffer_switch_done_latched_108 (.Q(buffer_switch_done_latched), 
           .C(SLM_CLK_c), .D(buffer_switch_done));   // src/usb3_if.v(70[8] 83[4])
    SB_LUT4 i1_2_lut_3_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[0]), 
            .I2(state_timeout_counter[2]), .I3(GND_net), .O(n4454));   // src/usb3_if.v(179[42:69])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h1e1e;
    SB_LUT4 sub_117_add_2_6_lut (.I0(GND_net), .I1(num_lines_clocked_out[4]), 
            .I2(VCC_net), .I3(n12115), .O(num_lines_clocked_out_10__N_441[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_117_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1565_2_lut_3_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[0]), 
            .I2(state_timeout_counter[2]), .I3(GND_net), .O(n6));   // src/usb3_if.v(179[42:69])
    defparam i1565_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY sub_117_add_2_6 (.CI(n12115), .I0(num_lines_clocked_out[4]), 
            .I1(VCC_net), .CO(n12116));
    SB_DFFSS state_FSM_i1 (.Q(n650[0]), .C(FIFO_CLK_c), .D(n3462), .S(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFESR dc32_fifo_data_in_latched__i31 (.Q(dc32_fifo_data_in_latched[31]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[31]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 sub_117_add_2_5_lut (.I0(GND_net), .I1(num_lines_clocked_out[3]), 
            .I2(VCC_net), .I3(n12114), .O(num_lines_clocked_out_10__N_441[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_117_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR dc32_fifo_data_in_latched__i30 (.Q(dc32_fifo_data_in_latched[30]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[30]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 mux_1382_i5_4_lut (.I0(n2737), .I1(state_timeout_counter[4]), 
            .I2(n2741), .I3(n8), .O(n2727));   // src/usb3_if.v(97[9] 199[16])
    defparam mux_1382_i5_4_lut.LUT_INIT = 16'hca3a;
    SB_LUT4 i7365_2_lut (.I0(n187[0]), .I1(n2744), .I2(GND_net), .I3(GND_net), 
            .O(n2737));   // src/usb3_if.v(173[26] 175[24])
    defparam i7365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_1382_i4_4_lut (.I0(n2737), .I1(state_timeout_counter[3]), 
            .I2(n2741), .I3(n6), .O(n2726));   // src/usb3_if.v(97[9] 199[16])
    defparam mux_1382_i4_4_lut.LUT_INIT = 16'hca3a;
    SB_LUT4 mux_1382_i3_4_lut (.I0(n2744), .I1(n4454), .I2(n2741), .I3(n187[0]), 
            .O(n2725));   // src/usb3_if.v(97[9] 199[16])
    defparam mux_1382_i3_4_lut.LUT_INIT = 16'h3f35;
    SB_DFFESR dc32_fifo_data_in_latched__i29 (.Q(dc32_fifo_data_in_latched[29]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[29]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i28 (.Q(dc32_fifo_data_in_latched[28]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[28]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i27 (.Q(dc32_fifo_data_in_latched[27]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[27]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i2083_3_lut (.I0(n609), .I1(DEBUG_1_c), .I2(n4226), .I3(GND_net), 
            .O(n2741));   // src/usb3_if.v(97[9] 199[16])
    defparam i2083_3_lut.LUT_INIT = 16'hbaba;
    SB_LUT4 i1_4_lut (.I0(n650[0]), .I1(n650[5]), .I2(n605), .I3(FT_OE_N_491), 
            .O(n12843));   // src/usb3_if.v(96[10] 200[8])
    defparam i1_4_lut.LUT_INIT = 16'h0ace;
    SB_LUT4 i4_4_lut (.I0(n650[8]), .I1(n663), .I2(n650[7]), .I3(reset_per_frame_latched), 
            .O(n10));   // src/usb3_if.v(96[10] 200[8])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12361_3_lut (.I0(n650[4]), .I1(n10), .I2(n12843), .I3(GND_net), 
            .O(n4839));   // src/usb3_if.v(96[10] 200[8])
    defparam i12361_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 mux_1382_i2_4_lut (.I0(n2744), .I1(state_timeout_counter[1]), 
            .I2(n2741), .I3(state_timeout_counter[0]), .O(n2724));   // src/usb3_if.v(97[9] 199[16])
    defparam mux_1382_i2_4_lut.LUT_INIT = 16'hca3a;
    SB_DFFESR dc32_fifo_data_in_latched__i26 (.Q(dc32_fifo_data_in_latched[26]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[26]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i25 (.Q(dc32_fifo_data_in_latched[25]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[25]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i24 (.Q(dc32_fifo_data_in_latched[24]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[24]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i23 (.Q(dc32_fifo_data_in_latched[23]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[23]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i22 (.Q(dc32_fifo_data_in_latched[22]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[22]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i21 (.Q(dc32_fifo_data_in_latched[21]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[21]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i20 (.Q(dc32_fifo_data_in_latched[20]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[20]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i19 (.Q(dc32_fifo_data_in_latched[19]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[19]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFSR write_to_dc32_fifo_latched_114 (.Q(write_to_dc32_fifo_latched), 
            .C(FIFO_CLK_c), .D(write_to_dc32_fifo_latched_N_503), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i18 (.Q(dc32_fifo_data_in_latched[18]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[18]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i17 (.Q(dc32_fifo_data_in_latched[17]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[17]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i16 (.Q(dc32_fifo_data_in_latched[16]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[16]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i15 (.Q(dc32_fifo_data_in_latched[15]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[15]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i14 (.Q(dc32_fifo_data_in_latched[14]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[14]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i13 (.Q(dc32_fifo_data_in_latched[13]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[13]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i12 (.Q(dc32_fifo_data_in_latched[12]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[12]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i11 (.Q(dc32_fifo_data_in_latched[11]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[11]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i10 (.Q(dc32_fifo_data_in_latched[10]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[10]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i9 (.Q(dc32_fifo_data_in_latched[9]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[9]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i8 (.Q(dc32_fifo_data_in_latched[8]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[8]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i7 (.Q(dc32_fifo_data_in_latched[7]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[7]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i6 (.Q(dc32_fifo_data_in_latched[6]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[6]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i5 (.Q(dc32_fifo_data_in_latched[5]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[5]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i4 (.Q(dc32_fifo_data_in_latched[4]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[4]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i3 (.Q(dc32_fifo_data_in_latched[3]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[3]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i2149_3_lut (.I0(n3611), .I1(n70[3]), .I2(n5298), .I3(GND_net), 
            .O(num_words_curr_line_5__N_435[3]));   // src/usb3_if.v(97[9] 199[16])
    defparam i2149_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR dc32_fifo_data_in_latched__i2 (.Q(dc32_fifo_data_in_latched[2]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[2]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i1 (.Q(dc32_fifo_data_in_latched[1]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[1]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i3951_3_lut (.I0(n4963), .I1(n5298), .I2(reset_per_frame_latched), 
            .I3(GND_net), .O(n5425));   // src/usb3_if.v(86[8] 201[4])
    defparam i3951_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 i3837_3_lut (.I0(FT_OE_N_495), .I1(n650[5]), .I2(n663), .I3(GND_net), 
            .O(n5298));   // src/usb3_if.v(97[9] 199[16])
    defparam i3837_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 i7443_3_lut (.I0(n172), .I1(n663), .I2(FT_OE_N_495), .I3(GND_net), 
            .O(n3611));   // src/usb3_if.v(97[9] 199[16])
    defparam i7443_3_lut.LUT_INIT = 16'hcdcd;
    SB_LUT4 i12222_4_lut (.I0(n172), .I1(n663), .I2(n12877), .I3(FT_OE_N_495), 
            .O(n14301));
    defparam i12222_4_lut.LUT_INIT = 16'hfcdc;
    SB_LUT4 i1_4_lut_adj_49 (.I0(reset_per_frame_latched), .I1(n14301), 
            .I2(FT_OE_N_491), .I3(n650[5]), .O(n4963));
    defparam i1_4_lut_adj_49.LUT_INIT = 16'hafee;
    SB_LUT4 i2153_3_lut (.I0(n3611), .I1(n70[5]), .I2(n5298), .I3(GND_net), 
            .O(num_words_curr_line_5__N_435[5]));   // src/usb3_if.v(97[9] 199[16])
    defparam i2153_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_117_add_2_5 (.CI(n12114), .I0(num_lines_clocked_out[3]), 
            .I1(VCC_net), .CO(n12115));
    SB_LUT4 sub_117_add_2_4_lut (.I0(GND_net), .I1(num_lines_clocked_out[2]), 
            .I2(VCC_net), .I3(n12113), .O(num_lines_clocked_out_10__N_441[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_117_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF state_FSM_i5 (.Q(n650[4]), .C(FIFO_CLK_c), .D(n7014));   // src/usb3_if.v(97[9] 199[16])
    SB_LUT4 i12312_2_lut_3_lut (.I0(num_words_curr_line[0]), .I1(n4772), 
            .I2(dc32_fifo_empty), .I3(GND_net), .O(n172));   // src/usb3_if.v(161[31:57])
    defparam i12312_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1932_3_lut_4_lut (.I0(num_words_curr_line[0]), .I1(n4772), 
            .I2(n650[2]), .I3(FR_RXF_c), .O(n4226));   // src/usb3_if.v(161[31:57])
    defparam i1932_3_lut_4_lut.LUT_INIT = 16'he0ef;
    SB_LUT4 FT_OE_I_8_2_lut_3_lut (.I0(num_words_curr_line[0]), .I1(n4772), 
            .I2(DEBUG_1_c), .I3(GND_net), .O(FT_OE_N_495));   // src/usb3_if.v(161[31:57])
    defparam FT_OE_I_8_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_CARRY sub_117_add_2_4 (.CI(n12113), .I0(num_lines_clocked_out[2]), 
            .I1(VCC_net), .CO(n12114));
    SB_LUT4 sub_117_add_2_3_lut (.I0(GND_net), .I1(num_lines_clocked_out[1]), 
            .I2(VCC_net), .I3(n12112), .O(num_lines_clocked_out_10__N_441[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_117_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_117_add_2_3 (.CI(n12112), .I0(num_lines_clocked_out[1]), 
            .I1(VCC_net), .CO(n12113));
    SB_LUT4 sub_117_add_2_2_lut (.I0(GND_net), .I1(num_lines_clocked_out[0]), 
            .I2(n172), .I3(VCC_net), .O(num_lines_clocked_out_10__N_441[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_117_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_117_add_2_2 (.CI(VCC_net), .I0(num_lines_clocked_out[0]), 
            .I1(n172), .CO(n12112));
    SB_LUT4 sub_114_add_2_7_lut (.I0(GND_net), .I1(num_words_curr_line[5]), 
            .I2(VCC_net), .I3(n12111), .O(n70[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_114_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_114_add_2_6_lut (.I0(GND_net), .I1(num_words_curr_line[4]), 
            .I2(VCC_net), .I3(n12110), .O(n70[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_114_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_114_add_2_6 (.CI(n12110), .I0(num_words_curr_line[4]), 
            .I1(VCC_net), .CO(n12111));
    SB_LUT4 sub_114_add_2_5_lut (.I0(GND_net), .I1(num_words_curr_line[3]), 
            .I2(VCC_net), .I3(n12109), .O(n70[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_114_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR num_lines_clocked_out_i10 (.Q(num_lines_clocked_out[10]), .C(FIFO_CLK_c), 
            .E(n4983), .D(num_lines_clocked_out_10__N_441[10]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i9 (.Q(num_lines_clocked_out[9]), .C(FIFO_CLK_c), 
            .E(n4983), .D(num_lines_clocked_out_10__N_441[9]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i8 (.Q(num_lines_clocked_out[8]), .C(FIFO_CLK_c), 
            .E(n4983), .D(num_lines_clocked_out_10__N_441[8]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i7 (.Q(num_lines_clocked_out[7]), .C(FIFO_CLK_c), 
            .E(n4983), .D(num_lines_clocked_out_10__N_441[7]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_CARRY sub_114_add_2_5 (.CI(n12109), .I0(num_words_curr_line[3]), 
            .I1(VCC_net), .CO(n12110));
    SB_DFFESR num_lines_clocked_out_i6 (.Q(num_lines_clocked_out[6]), .C(FIFO_CLK_c), 
            .E(n4983), .D(num_lines_clocked_out_10__N_441[6]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 sub_114_add_2_4_lut (.I0(GND_net), .I1(num_words_curr_line[2]), 
            .I2(VCC_net), .I3(n12108), .O(n70[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_114_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS num_lines_clocked_out_i5 (.Q(num_lines_clocked_out[5]), .C(FIFO_CLK_c), 
            .E(n4983), .D(num_lines_clocked_out_10__N_441[5]), .S(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i4 (.Q(num_lines_clocked_out[4]), .C(FIFO_CLK_c), 
            .E(n4983), .D(num_lines_clocked_out_10__N_441[4]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i3 (.Q(num_lines_clocked_out[3]), .C(FIFO_CLK_c), 
            .E(n4983), .D(num_lines_clocked_out_10__N_441[3]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i2 (.Q(num_lines_clocked_out[2]), .C(FIFO_CLK_c), 
            .E(n4983), .D(num_lines_clocked_out_10__N_441[2]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i1 (.Q(num_lines_clocked_out[1]), .C(FIFO_CLK_c), 
            .E(n4983), .D(num_lines_clocked_out_10__N_441[1]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESS num_words_curr_line_i5 (.Q(num_words_curr_line[5]), .C(FIFO_CLK_c), 
            .E(n4963), .D(num_words_curr_line_5__N_435[5]), .S(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_words_curr_line_i4 (.Q(num_words_curr_line[4]), .C(FIFO_CLK_c), 
            .E(n4963), .D(n70[4]), .R(n5425));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESS num_words_curr_line_i3 (.Q(num_words_curr_line[3]), .C(FIFO_CLK_c), 
            .E(n4963), .D(num_words_curr_line_5__N_435[3]), .S(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_words_curr_line_i2 (.Q(num_words_curr_line[2]), .C(FIFO_CLK_c), 
            .E(n4963), .D(n70[2]), .R(n5425));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_words_curr_line_i1 (.Q(num_words_curr_line[1]), .C(FIFO_CLK_c), 
            .E(n4963), .D(n70[1]), .R(n5425));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i245_4_lut (.I0(n8999), .I1(n11), .I2(n650[5]), .I3(FR_RXF_c), 
            .O(write_to_dc32_fifo_latched_N_503));   // src/usb3_if.v(97[9] 199[16])
    defparam i245_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY sub_114_add_2_4 (.CI(n12108), .I0(num_words_curr_line[2]), 
            .I1(VCC_net), .CO(n12109));
    SB_LUT4 sub_114_add_2_3_lut (.I0(GND_net), .I1(num_words_curr_line[1]), 
            .I2(VCC_net), .I3(n12107), .O(n70[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_114_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(FIFO_CLK_c), 
            .E(n4839), .D(n2724), .R(n5368));   // src/usb3_if.v(86[8] 201[4])
    SB_CARRY sub_114_add_2_3 (.CI(n12107), .I0(num_words_curr_line[1]), 
            .I1(VCC_net), .CO(n12108));
    SB_LUT4 sub_114_add_2_2_lut (.I0(GND_net), .I1(num_words_curr_line[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n70[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_114_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_114_add_2_2 (.CI(VCC_net), .I0(num_words_curr_line[0]), 
            .I1(GND_net), .CO(n12107));
    SB_DFFESS state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(FIFO_CLK_c), 
            .E(n4839), .D(n2725), .S(n5368));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(FIFO_CLK_c), 
            .E(n4839), .D(n2726), .R(n5368));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(FIFO_CLK_c), 
            .E(n4839), .D(n2727), .R(n5368));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i0 (.Q(dc32_fifo_data_in_latched[0]), 
            .C(FIFO_CLK_c), .E(n5138), .D(n850[0]), .R(n5387));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i2_3_lut (.I0(n650[5]), .I1(n650[6]), .I2(n650[4]), .I3(GND_net), 
            .O(n883));   // src/usb3_if.v(97[9] 199[16])
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3913_3_lut (.I0(n5138), .I1(n883), .I2(reset_per_frame_latched), 
            .I3(GND_net), .O(n5387));   // src/usb3_if.v(86[8] 201[4])
    defparam i3913_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 i2_3_lut_adj_50 (.I0(reset_per_frame_latched), .I1(n650[2]), 
            .I2(n883), .I3(GND_net), .O(n5138));
    defparam i2_3_lut_adj_50.LUT_INIT = 16'hfbfb;
    SB_LUT4 i7_4_lut (.I0(num_lines_clocked_out[7]), .I1(num_lines_clocked_out[2]), 
            .I2(num_lines_clocked_out[9]), .I3(num_lines_clocked_out[0]), 
            .O(n18));   // src/usb3_if.v(164[29:57])
    defparam i7_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i5_2_lut (.I0(num_lines_clocked_out[1]), .I1(num_lines_clocked_out[5]), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // src/usb3_if.v(164[29:57])
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut (.I0(num_lines_clocked_out[6]), .I1(n18), .I2(num_lines_clocked_out[3]), 
            .I3(num_lines_clocked_out[10]), .O(n20));   // src/usb3_if.v(164[29:57])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(num_lines_clocked_out[4]), .I1(n20), .I2(n16), 
            .I3(num_lines_clocked_out[8]), .O(n187[0]));   // src/usb3_if.v(164[29:57])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2011_4_lut (.I0(n650[0]), .I1(n187[0]), .I2(n607), .I3(n2744), 
            .O(n3462));   // src/usb3_if.v(97[9] 199[16])
    defparam i2011_4_lut.LUT_INIT = 16'hb3a0;
    SB_DFFN dc32_fifo_data_in_i1 (.Q(dc32_fifo_data_in[1]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[1]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i2 (.Q(dc32_fifo_data_in[2]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[2]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i3 (.Q(dc32_fifo_data_in[3]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[3]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i4 (.Q(dc32_fifo_data_in[4]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[4]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i5 (.Q(dc32_fifo_data_in[5]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[5]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i6 (.Q(dc32_fifo_data_in[6]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[6]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i7 (.Q(dc32_fifo_data_in[7]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[7]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i8 (.Q(dc32_fifo_data_in[8]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[8]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i9 (.Q(dc32_fifo_data_in[9]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[9]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i10 (.Q(dc32_fifo_data_in[10]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[10]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i11 (.Q(dc32_fifo_data_in[11]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[11]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i12 (.Q(dc32_fifo_data_in[12]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[12]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i13 (.Q(dc32_fifo_data_in[13]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[13]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i14 (.Q(dc32_fifo_data_in[14]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[14]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i15 (.Q(dc32_fifo_data_in[15]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[15]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i16 (.Q(dc32_fifo_data_in[16]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[16]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i17 (.Q(dc32_fifo_data_in[17]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[17]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i18 (.Q(dc32_fifo_data_in[18]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[18]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i19 (.Q(dc32_fifo_data_in[19]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[19]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i20 (.Q(dc32_fifo_data_in[20]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[20]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i21 (.Q(dc32_fifo_data_in[21]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[21]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i22 (.Q(dc32_fifo_data_in[22]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[22]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i23 (.Q(dc32_fifo_data_in[23]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[23]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i24 (.Q(dc32_fifo_data_in[24]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[24]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i25 (.Q(dc32_fifo_data_in[25]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[25]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i26 (.Q(dc32_fifo_data_in[26]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[26]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i27 (.Q(dc32_fifo_data_in[27]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[27]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i28 (.Q(dc32_fifo_data_in[28]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[28]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i29 (.Q(dc32_fifo_data_in[29]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[29]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i30 (.Q(dc32_fifo_data_in[30]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[30]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i31 (.Q(dc32_fifo_data_in[31]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[31]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFESS FT_OE_111 (.Q(FT_OE_c), .C(FIFO_CLK_c), .E(VCC_net), .D(FT_OE_N_490), 
            .S(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 sub_117_add_2_12_lut (.I0(GND_net), .I1(num_lines_clocked_out[10]), 
            .I2(VCC_net), .I3(n12121), .O(num_lines_clocked_out_10__N_441[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_117_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR num_lines_clocked_out_i0 (.Q(num_lines_clocked_out[0]), .C(FIFO_CLK_c), 
            .E(n4983), .D(num_lines_clocked_out_10__N_441[0]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_words_curr_line_i0 (.Q(num_words_curr_line[0]), .C(FIFO_CLK_c), 
            .E(n4963), .D(n70[0]), .R(n5425));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 sub_117_add_2_11_lut (.I0(GND_net), .I1(num_lines_clocked_out[9]), 
            .I2(VCC_net), .I3(n12120), .O(num_lines_clocked_out_10__N_441[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_117_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_117_add_2_11 (.CI(n12120), .I0(num_lines_clocked_out[9]), 
            .I1(VCC_net), .CO(n12121));
    SB_LUT4 sub_117_add_2_10_lut (.I0(GND_net), .I1(num_lines_clocked_out[8]), 
            .I2(VCC_net), .I3(n12119), .O(num_lines_clocked_out_10__N_441[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_117_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(FIFO_CLK_c), 
            .E(n4839), .D(n2723), .R(n5368));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFSR state_FSM_i2 (.Q(n650[1]), .C(FIFO_CLK_c), .D(n12840), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFSR state_FSM_i3 (.Q(n650[2]), .C(FIFO_CLK_c), .D(n3458), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFSR state_FSM_i4 (.Q(n663), .C(FIFO_CLK_c), .D(n696), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFSR state_FSM_i6 (.Q(n650[5]), .C(FIFO_CLK_c), .D(n3456), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFSR state_FSM_i7 (.Q(n650[6]), .C(FIFO_CLK_c), .D(n3452), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFSR state_FSM_i8 (.Q(n650[7]), .C(FIFO_CLK_c), .D(n706), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFSR state_FSM_i9 (.Q(n650[8]), .C(FIFO_CLK_c), .D(n709), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_LUT4 i158_2_lut_3_lut (.I0(buffer_switch_done_latched), .I1(dc32_fifo_empty_latched), 
            .I2(FR_RXF_c), .I3(GND_net), .O(n607));   // src/usb3_if.v(99[21:96])
    defparam i158_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i156_2_lut_3_lut (.I0(buffer_switch_done_latched), .I1(dc32_fifo_empty_latched), 
            .I2(FR_RXF_c), .I3(GND_net), .O(n605));   // src/usb3_if.v(99[21:96])
    defparam i156_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_1361));   // src/usb3_if.v(153[21:49])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_51 (.I0(state_timeout_counter[3]), .I1(state_timeout_counter[2]), 
            .I2(state_timeout_counter[0]), .I3(n6_adj_1361), .O(n609));   // src/usb3_if.v(153[21:49])
    defparam i4_4_lut_adj_51.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_adj_52 (.I0(n650[2]), .I1(n609), .I2(GND_net), .I3(GND_net), 
            .O(n12877));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_2_lut_adj_52.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_53 (.I0(num_words_curr_line[5]), .I1(num_words_curr_line[1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_1362));   // src/usb3_if.v(161[31:57])
    defparam i1_2_lut_adj_53.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_54 (.I0(num_words_curr_line[3]), .I1(num_words_curr_line[4]), 
            .I2(num_words_curr_line[2]), .I3(n6_adj_1362), .O(n4772));   // src/usb3_if.v(161[31:57])
    defparam i4_4_lut_adj_54.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_55 (.I0(num_words_curr_line[0]), .I1(n4772), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // src/usb3_if.v(132[21:47])
    defparam i1_2_lut_adj_55.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_56 (.I0(n650[4]), .I1(n650[8]), .I2(GND_net), 
            .I3(GND_net), .O(n918));
    defparam i1_2_lut_adj_56.LUT_INIT = 16'heeee;
    SB_LUT4 i7522_2_lut_3_lut (.I0(FT_OE_N_495), .I1(n609), .I2(n172), 
            .I3(GND_net), .O(n8991));   // src/usb3_if.v(153[17] 176[20])
    defparam i7522_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_3_lut_4_lut (.I0(FT_OE_N_495), .I1(n609), .I2(n650[2]), 
            .I3(reset_per_frame_latched), .O(n4983));   // src/usb3_if.v(153[17] 176[20])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hff10;
    SB_LUT4 i2_3_lut_4_lut (.I0(FT_OE_N_495), .I1(n609), .I2(n172), .I3(n650[2]), 
            .O(n2744));   // src/usb3_if.v(153[17] 176[20])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1956_4_lut (.I0(n8999), .I1(FT_OE_N_491), .I2(n650[5]), .I3(n918), 
            .O(FT_RD_N_501));   // src/usb3_if.v(97[9] 199[16])
    defparam i1956_4_lut.LUT_INIT = 16'hc0c5;
    SB_CARRY sub_117_add_2_10 (.CI(n12119), .I0(num_lines_clocked_out[8]), 
            .I1(VCC_net), .CO(n12120));
    SB_LUT4 sub_117_add_2_9_lut (.I0(GND_net), .I1(num_lines_clocked_out[7]), 
            .I2(VCC_net), .I3(n12118), .O(num_lines_clocked_out_10__N_441[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_117_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_117_add_2_9 (.CI(n12118), .I0(num_lines_clocked_out[7]), 
            .I1(VCC_net), .CO(n12119));
    SB_LUT4 sub_117_add_2_8_lut (.I0(GND_net), .I1(num_lines_clocked_out[6]), 
            .I2(VCC_net), .I3(n12117), .O(num_lines_clocked_out_10__N_441[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_117_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_117_add_2_8 (.CI(n12117), .I0(num_lines_clocked_out[6]), 
            .I1(VCC_net), .CO(n12118));
    SB_LUT4 sub_117_add_2_7_lut (.I0(GND_net), .I1(num_lines_clocked_out[5]), 
            .I2(VCC_net), .I3(n12116), .O(num_lines_clocked_out_10__N_441[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_117_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7196_2_lut_3_lut_4_lut (.I0(DEBUG_3_c_0_c), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[0]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7196_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7332_2_lut_3_lut_4_lut (.I0(FIFO_D1_c_1), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[1]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7332_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7333_2_lut_3_lut_4_lut (.I0(FIFO_D2_c_2), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[2]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7333_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7334_2_lut_3_lut_4_lut (.I0(FIFO_D3_c_3), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[3]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7334_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7335_2_lut_3_lut_4_lut (.I0(FIFO_D4_c_4), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[4]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7335_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7336_2_lut_3_lut_4_lut (.I0(FIFO_D5_c_5), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[5]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7336_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7337_2_lut_3_lut_4_lut (.I0(FIFO_D6_c_6), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[6]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7337_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7338_2_lut_3_lut_4_lut (.I0(FIFO_D7_c_7), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[7]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7338_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7339_2_lut_3_lut_4_lut (.I0(FIFO_D8_c_8), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[8]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7339_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_CARRY sub_117_add_2_7 (.CI(n12116), .I0(num_lines_clocked_out[5]), 
            .I1(VCC_net), .CO(n12117));
    SB_LUT4 i7340_2_lut_3_lut_4_lut (.I0(FIFO_D9_c_9), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[9]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7340_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7341_2_lut_3_lut_4_lut (.I0(FIFO_D10_c_10), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[10]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7341_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7342_2_lut_3_lut_4_lut (.I0(FIFO_D11_c_11), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[11]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7342_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7343_2_lut_3_lut_4_lut (.I0(FIFO_D12_c_12), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[12]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7343_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7344_2_lut_3_lut_4_lut (.I0(FIFO_D13_c_13), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[13]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7344_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7345_2_lut_3_lut_4_lut (.I0(FIFO_D14_c_14), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[14]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7345_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7346_2_lut_3_lut_4_lut (.I0(FIFO_D15_c_15), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[15]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7346_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7347_2_lut_3_lut_4_lut (.I0(FIFO_D16_c_16), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[16]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7347_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7348_2_lut_3_lut_4_lut (.I0(FIFO_D17_c_17), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[17]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7348_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7349_2_lut_3_lut_4_lut (.I0(FIFO_D18_c_18), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[18]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7349_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7350_2_lut_3_lut_4_lut (.I0(FIFO_D19_c_19), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[19]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7350_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7351_2_lut_3_lut_4_lut (.I0(FIFO_D20_c_20), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[20]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7351_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7352_2_lut_3_lut_4_lut (.I0(FIFO_D21_c_21), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[21]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7352_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7353_2_lut_3_lut_4_lut (.I0(FIFO_D22_c_22), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[22]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7353_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7354_2_lut_3_lut_4_lut (.I0(FIFO_D23_c_23), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[23]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7354_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7355_2_lut_3_lut_4_lut (.I0(FIFO_D24_c_24), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[24]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7355_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7356_2_lut_3_lut_4_lut (.I0(FIFO_D25_c_25), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[25]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7356_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i1_2_lut_3_lut_adj_57 (.I0(n650[5]), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(GND_net), .O(n4757));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_2_lut_3_lut_adj_57.LUT_INIT = 16'ha2a2;
    SB_LUT4 i2005_3_lut_4_lut (.I0(FR_RXF_c), .I1(n650[4]), .I2(n650[8]), 
            .I3(n4757), .O(n3456));   // src/usb3_if.v(97[9] 199[16])
    defparam i2005_3_lut_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i7357_2_lut_3_lut_4_lut (.I0(FIFO_D26_c_26), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[26]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7357_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i263_4_lut (.I0(FT_OE_N_491), .I1(n8999), .I2(n12270), .I3(n650[5]), 
            .O(FT_OE_N_490));   // src/usb3_if.v(97[9] 199[16])
    defparam i263_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i7358_2_lut_3_lut_4_lut (.I0(FIFO_D27_c_27), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[27]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7358_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7359_2_lut_3_lut_4_lut (.I0(FIFO_D28_c_28), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[28]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7359_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7360_2_lut_3_lut_4_lut (.I0(FIFO_D29_c_29), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[29]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7360_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i7361_2_lut_3_lut_4_lut (.I0(FIFO_D30_c_30), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[30]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7361_2_lut_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i1_2_lut_3_lut_adj_58 (.I0(FT_OE_N_495), .I1(n650[2]), .I2(n609), 
            .I3(GND_net), .O(n8999));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_2_lut_3_lut_adj_58.LUT_INIT = 16'h0808;
    SB_LUT4 i7197_2_lut_3_lut (.I0(FR_RXF_c), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(GND_net), .O(FT_OE_N_491));   // src/usb3_if.v(137[22] 148[20])
    defparam i7197_2_lut_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i7362_2_lut_4_lut (.I0(FIFO_D31_c_31), .I1(num_words_curr_line[0]), 
            .I2(n4772), .I3(n650[5]), .O(n850[31]));   // src/usb3_if.v(137[22] 148[20])
    defparam i7362_2_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i211_2_lut_3_lut (.I0(num_words_curr_line[0]), .I1(n4772), .I2(n650[5]), 
            .I3(GND_net), .O(n694));   // src/usb3_if.v(97[9] 199[16])
    defparam i211_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 mux_1382_i1_3_lut (.I0(n2744), .I1(state_timeout_counter[0]), 
            .I2(n2741), .I3(GND_net), .O(n2723));   // src/usb3_if.v(97[9] 199[16])
    defparam mux_1382_i1_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_4_lut_adj_59 (.I0(n2737), .I1(n605), .I2(n3459), .I3(n650[0]), 
            .O(n12840));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_4_lut_adj_59.LUT_INIT = 16'hfefa;
    SB_LUT4 i2008_2_lut (.I0(n650[1]), .I1(n8685), .I2(GND_net), .I3(GND_net), 
            .O(n3459));   // src/usb3_if.v(97[9] 199[16])
    defparam i2008_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7219_3_lut (.I0(FR_RXF_c), .I1(n609), .I2(DEBUG_1_c), .I3(GND_net), 
            .O(n8685));
    defparam i7219_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2007_4_lut (.I0(n650[2]), .I1(n694), .I2(n609), .I3(n8991), 
            .O(n3458));   // src/usb3_if.v(97[9] 199[16])
    defparam i2007_4_lut.LUT_INIT = 16'hecee;
    SB_LUT4 i213_2_lut (.I0(n8685), .I1(n650[1]), .I2(GND_net), .I3(GND_net), 
            .O(n696));   // src/usb3_if.v(97[9] 199[16])
    defparam i213_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2001_4_lut (.I0(n650[6]), .I1(FR_RXF_c), .I2(n8685), .I3(n4757), 
            .O(n3452));   // src/usb3_if.v(97[9] 199[16])
    defparam i2001_4_lut.LUT_INIT = 16'heca0;
    SB_LUT4 i223_2_lut (.I0(n8685), .I1(n650[6]), .I2(GND_net), .I3(GND_net), 
            .O(n706));   // src/usb3_if.v(97[9] 199[16])
    defparam i223_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 reduce_or_225_i1_2_lut (.I0(n650[7]), .I1(n8999), .I2(GND_net), 
            .I3(GND_net), .O(n709));   // src/usb3_if.v(97[9] 199[16])
    defparam reduce_or_225_i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_4_lut_adj_60 (.I0(n650[0]), .I1(n650[2]), .I2(n650[1]), 
            .I3(n650[6]), .O(n12270));
    defparam i2_3_lut_4_lut_adj_60.LUT_INIT = 16'hfffe;
    SB_LUT4 i1573_2_lut_4_lut (.I0(state_timeout_counter[3]), .I1(state_timeout_counter[1]), 
            .I2(state_timeout_counter[0]), .I3(state_timeout_counter[2]), 
            .O(n8));   // src/usb3_if.v(179[42:69])
    defparam i1573_2_lut_4_lut.LUT_INIT = 16'hfffe;
    
endmodule
//
// Verilog Description of module clock
//

module clock (GND_net, VCC_net, ICE_SYSCLK_c, pll_clk_unbuf) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    input ICE_SYSCLK_c;
    output pll_clk_unbuf;
    
    
    SB_PLL40_CORE pll_config (.REFERENCECLK(ICE_SYSCLK_c), .PLLOUTGLOBAL(pll_clk_unbuf), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=15, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=222, LSE_RLINE=228 */ ;   // src/top.v(222[7] 228[3])
    defparam pll_config.FEEDBACK_PATH = "SIMPLE";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll_config.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll_config.FDA_FEEDBACK = 0;
    defparam pll_config.FDA_RELATIVE = 0;
    defparam pll_config.PLLOUT_SELECT = "GENCLK";
    defparam pll_config.DIVR = 4'b0001;
    defparam pll_config.DIVF = 7'b1010010;
    defparam pll_config.DIVQ = 3'b100;
    defparam pll_config.FILTER_RANGE = 3'b001;
    defparam pll_config.ENABLE_ICEGATE = 1'b0;
    defparam pll_config.TEST_MODE = 1'b0;
    defparam pll_config.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module spi
//

module spi (n4837, SLM_CLK_c, GND_net, tx_addr_byte, n2407, SEN_c_1, 
            \tx_data_byte[7] , SOUT_c, n4884, \rx_shift_reg[0] , SDAT_c_15, 
            n6988, rx_buf_byte, n6987, n6986, n6985, n6984, n6983, 
            n6982, n6981, \rx_shift_reg[7] , n6980, \rx_shift_reg[6] , 
            n6979, \rx_shift_reg[5] , n6978, \rx_shift_reg[4] , n6977, 
            \rx_shift_reg[3] , n6976, \rx_shift_reg[2] , n6975, \rx_shift_reg[1] , 
            n12537, VCC_net, \tx_shift_reg[0] , \tx_data_byte[1] , multi_byte_spi_trans_flag_r, 
            \tx_data_byte[2] , \tx_data_byte[3] , \tx_data_byte[4] , spi_rx_byte_ready, 
            SCK_c_0, spi_start_transfer_r, n5578, \tx_data_byte[5] , 
            \tx_data_byte[6] , n3963) /* synthesis syn_module_defined=1 */ ;
    output n4837;
    input SLM_CLK_c;
    input GND_net;
    input [7:0]tx_addr_byte;
    output n2407;
    output SEN_c_1;
    input \tx_data_byte[7] ;
    input SOUT_c;
    output n4884;
    output \rx_shift_reg[0] ;
    output SDAT_c_15;
    input n6988;
    output [7:0]rx_buf_byte;
    input n6987;
    input n6986;
    input n6985;
    input n6984;
    input n6983;
    input n6982;
    input n6981;
    output \rx_shift_reg[7] ;
    input n6980;
    output \rx_shift_reg[6] ;
    input n6979;
    output \rx_shift_reg[5] ;
    input n6978;
    output \rx_shift_reg[4] ;
    input n6977;
    output \rx_shift_reg[3] ;
    input n6976;
    output \rx_shift_reg[2] ;
    input n6975;
    output \rx_shift_reg[1] ;
    input n12537;
    input VCC_net;
    output \tx_shift_reg[0] ;
    input \tx_data_byte[1] ;
    input multi_byte_spi_trans_flag_r;
    input \tx_data_byte[2] ;
    input \tx_data_byte[3] ;
    input \tx_data_byte[4] ;
    output spi_rx_byte_ready;
    output SCK_c_0;
    input spi_start_transfer_r;
    input n5578;
    input \tx_data_byte[5] ;
    input \tx_data_byte[6] ;
    output n3963;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [15:0]n2408;
    wire [15:0]tx_shift_reg;   // src/spi.v(70[12:24])
    wire [3:0]state;   // src/spi.v(71[11:16])
    
    wire n14, n19, n14252, n14253, n34;
    wire [7:0]n2484;
    
    wire n37, n12966, n5394, n4776, n4912;
    wire [2:0]n1140;
    wire [3:0]state_3__N_1123;
    
    wire n16230, n5054, n5383, n14300;
    wire [7:0]n315;
    wire [7:0]multi_byte_counter;   // src/spi.v(68[11:29])
    
    wire n12143, n12142;
    wire [9:0]n45;
    wire [9:0]counter;   // src/spi.v(69[11:18])
    
    wire n12186, n12185, n3, n3_adj_1353, n21, n12184, n12141, 
        n12183, n12182, n12140, n12139, n12181, n12180, n12179, 
        n12138, n12178, n12137, n12890, n12889, n19_adj_1354, n13000, 
        n12820, n13004, n4896, n6, n5062, n12829, n4570, n4705, 
        n10, n14_adj_1355, n10_adj_1356, n14_adj_1357, n14298, n7, 
        n14305, n24, n4, n16, n24_adj_1358, n8, n14272, n13036, 
        n7_adj_1359, n14309, n12888, n3_adj_1360, n22, n14271;
    
    SB_DFFE tx_shift_reg_i0_i6 (.Q(tx_shift_reg[6]), .C(SLM_CLK_c), .E(n4837), 
            .D(n2408[6]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i5 (.Q(tx_shift_reg[5]), .C(SLM_CLK_c), .E(n4837), 
            .D(n2408[5]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i1_3_lut (.I0(state[3]), .I1(state[2]), .I2(state[0]), .I3(GND_net), 
            .O(n14));   // src/spi.v(88[9] 219[16])
    defparam i1_3_lut.LUT_INIT = 16'hcdcd;
    SB_LUT4 i12217_3_lut (.I0(state[0]), .I1(state[2]), .I2(n19), .I3(GND_net), 
            .O(n14252));
    defparam i12217_3_lut.LUT_INIT = 16'h4d4d;
    SB_LUT4 i12218_3_lut (.I0(state[3]), .I1(state[2]), .I2(state[0]), 
            .I3(GND_net), .O(n14253));
    defparam i12218_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i65_3_lut (.I0(n14), .I1(n14252), .I2(state[1]), .I3(GND_net), 
            .O(n34));
    defparam i65_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i66_4_lut (.I0(n14253), .I1(n2484[4]), .I2(state[1]), .I3(state[3]), 
            .O(n37));
    defparam i66_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_4_lut (.I0(state[3]), .I1(n37), .I2(n34), .I3(n12966), 
            .O(n5394));
    defparam i1_4_lut.LUT_INIT = 16'h50dc;
    SB_LUT4 i12332_4_lut (.I0(state[3]), .I1(state[1]), .I2(n4776), .I3(n14), 
            .O(n4912));   // src/spi.v(88[9] 219[16])
    defparam i12332_4_lut.LUT_INIT = 16'h4c5f;
    SB_LUT4 mux_1164_i15_3_lut (.I0(tx_addr_byte[6]), .I1(tx_shift_reg[13]), 
            .I2(n2407), .I3(GND_net), .O(n2408[14]));   // src/spi.v(88[9] 219[16])
    defparam mux_1164_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1164_i14_3_lut (.I0(tx_addr_byte[5]), .I1(tx_shift_reg[12]), 
            .I2(n2407), .I3(GND_net), .O(n2408[13]));   // src/spi.v(88[9] 219[16])
    defparam mux_1164_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1164_i13_3_lut (.I0(tx_addr_byte[4]), .I1(tx_shift_reg[11]), 
            .I2(n2407), .I3(GND_net), .O(n2408[12]));   // src/spi.v(88[9] 219[16])
    defparam mux_1164_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1164_i12_3_lut (.I0(tx_addr_byte[3]), .I1(tx_shift_reg[10]), 
            .I2(n2407), .I3(GND_net), .O(n2408[11]));   // src/spi.v(88[9] 219[16])
    defparam mux_1164_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1164_i11_3_lut (.I0(tx_addr_byte[2]), .I1(tx_shift_reg[9]), 
            .I2(n2407), .I3(GND_net), .O(n2408[10]));   // src/spi.v(88[9] 219[16])
    defparam mux_1164_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1164_i10_3_lut (.I0(tx_addr_byte[1]), .I1(tx_shift_reg[8]), 
            .I2(n2407), .I3(GND_net), .O(n2408[9]));   // src/spi.v(88[9] 219[16])
    defparam mux_1164_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1164_i9_3_lut (.I0(tx_addr_byte[0]), .I1(tx_shift_reg[7]), 
            .I2(n2407), .I3(GND_net), .O(n2408[8]));   // src/spi.v(88[9] 219[16])
    defparam mux_1164_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF byte_recv_92_i2 (.Q(SEN_c_1), .C(SLM_CLK_c), .D(n1140[1]));   // src/spi.v(88[9] 219[16])
    SB_LUT4 mux_1164_i8_3_lut (.I0(\tx_data_byte[7] ), .I1(tx_shift_reg[6]), 
            .I2(n2407), .I3(GND_net), .O(n2408[7]));   // src/spi.v(88[9] 219[16])
    defparam mux_1164_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE rx_shift_reg_i0 (.Q(\rx_shift_reg[0] ), .C(SLM_CLK_c), .E(n4884), 
            .D(SOUT_c));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i0 (.Q(state[0]), .C(SLM_CLK_c), .E(n16230), .D(state_3__N_1123[0]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i4 (.Q(tx_shift_reg[4]), .C(SLM_CLK_c), .E(n4837), 
            .D(n2408[4]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i3 (.Q(tx_shift_reg[3]), .C(SLM_CLK_c), .E(n4837), 
            .D(n2408[3]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i2 (.Q(tx_shift_reg[2]), .C(SLM_CLK_c), .E(n4837), 
            .D(n2408[2]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i15 (.Q(SDAT_c_15), .C(SLM_CLK_c), .E(n4837), 
            .D(n2408[15]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i1 (.Q(tx_shift_reg[1]), .C(SLM_CLK_c), .E(n4837), 
            .D(n2408[1]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i10859_2_lut (.I0(state[0]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n12966));
    defparam i10859_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3909_2_lut (.I0(n5054), .I1(state[3]), .I2(GND_net), .I3(GND_net), 
            .O(n5383));   // src/spi.v(76[8] 221[4])
    defparam i3909_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_36 (.I0(state[1]), .I1(n14300), .I2(n12966), 
            .I3(state[3]), .O(n5054));
    defparam i1_4_lut_adj_36.LUT_INIT = 16'h0a88;
    SB_DFF Rx_Recv_Byte_i7 (.Q(rx_buf_byte[7]), .C(SLM_CLK_c), .D(n6988));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i6 (.Q(rx_buf_byte[6]), .C(SLM_CLK_c), .D(n6987));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i5 (.Q(rx_buf_byte[5]), .C(SLM_CLK_c), .D(n6986));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i4 (.Q(rx_buf_byte[4]), .C(SLM_CLK_c), .D(n6985));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i3 (.Q(rx_buf_byte[3]), .C(SLM_CLK_c), .D(n6984));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i2 (.Q(rx_buf_byte[2]), .C(SLM_CLK_c), .D(n6983));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i1 (.Q(rx_buf_byte[1]), .C(SLM_CLK_c), .D(n6982));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i7 (.Q(\rx_shift_reg[7] ), .C(SLM_CLK_c), .D(n6981));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i6 (.Q(\rx_shift_reg[6] ), .C(SLM_CLK_c), .D(n6980));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i5 (.Q(\rx_shift_reg[5] ), .C(SLM_CLK_c), .D(n6979));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i4 (.Q(\rx_shift_reg[4] ), .C(SLM_CLK_c), .D(n6978));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i3 (.Q(\rx_shift_reg[3] ), .C(SLM_CLK_c), .D(n6977));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i2 (.Q(\rx_shift_reg[2] ), .C(SLM_CLK_c), .D(n6976));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i1 (.Q(\rx_shift_reg[1] ), .C(SLM_CLK_c), .D(n6975));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i0 (.Q(\tx_shift_reg[0] ), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n12537));   // src/spi.v(76[8] 221[4])
    SB_DFFESS multi_byte_counter_i7 (.Q(multi_byte_counter[7]), .C(SLM_CLK_c), 
            .E(n5054), .D(n315[7]), .S(n5383));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i6 (.Q(multi_byte_counter[6]), .C(SLM_CLK_c), 
            .E(n5054), .D(n315[6]), .R(n5383));   // src/spi.v(76[8] 221[4])
    SB_DFFESS multi_byte_counter_i5 (.Q(multi_byte_counter[5]), .C(SLM_CLK_c), 
            .E(n5054), .D(n315[5]), .S(n5383));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i4 (.Q(multi_byte_counter[4]), .C(SLM_CLK_c), 
            .E(n5054), .D(n315[4]), .R(n5383));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i3 (.Q(multi_byte_counter[3]), .C(SLM_CLK_c), 
            .E(n5054), .D(n315[3]), .R(n5383));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i2 (.Q(multi_byte_counter[2]), .C(SLM_CLK_c), 
            .E(n5054), .D(n315[2]), .R(n5383));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i1 (.Q(multi_byte_counter[1]), .C(SLM_CLK_c), 
            .E(n5054), .D(n315[1]), .R(n5383));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_1164_i2_3_lut (.I0(\tx_data_byte[1] ), .I1(\tx_shift_reg[0] ), 
            .I2(n2407), .I3(GND_net), .O(n2408[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_1164_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1186_9_lut (.I0(GND_net), .I1(multi_byte_counter[7]), .I2(n2484[4]), 
            .I3(n12143), .O(n315[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1186_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1186_8_lut (.I0(GND_net), .I1(multi_byte_counter[6]), .I2(n2484[4]), 
            .I3(n12142), .O(n315[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1186_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1437_add_4_11_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[9]), 
            .I3(n12186), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1437_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1437_add_4_10_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[8]), 
            .I3(n12185), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1437_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_56_Mux_1_i3_3_lut_3_lut (.I0(multi_byte_spi_trans_flag_r), 
            .I1(state[0]), .I2(state[1]), .I3(GND_net), .O(n3));
    defparam mux_56_Mux_1_i3_3_lut_3_lut.LUT_INIT = 16'h3e3e;
    SB_CARRY add_1186_8 (.CI(n12142), .I0(multi_byte_counter[6]), .I1(n2484[4]), 
            .CO(n12143));
    SB_LUT4 mux_56_Mux_0_i3_4_lut_4_lut (.I0(multi_byte_spi_trans_flag_r), 
            .I1(state[0]), .I2(state[1]), .I3(n19), .O(n3_adj_1353));
    defparam mux_56_Mux_0_i3_4_lut_4_lut.LUT_INIT = 16'hc131;
    SB_CARRY counter_1437_add_4_10 (.CI(n12185), .I0(VCC_net), .I1(counter[8]), 
            .CO(n12186));
    SB_LUT4 i43_4_lut_4_lut (.I0(state[3]), .I1(state[2]), .I2(state[1]), 
            .I3(state[0]), .O(n21));
    defparam i43_4_lut_4_lut.LUT_INIT = 16'hf01a;
    SB_LUT4 counter_1437_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[7]), 
            .I3(n12184), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1437_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1186_7_lut (.I0(GND_net), .I1(multi_byte_counter[5]), .I2(n2484[4]), 
            .I3(n12141), .O(n315[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1186_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1437_add_4_9 (.CI(n12184), .I0(VCC_net), .I1(counter[7]), 
            .CO(n12185));
    SB_LUT4 counter_1437_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[6]), 
            .I3(n12183), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1437_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3861_3_lut_4_lut (.I0(state[3]), .I1(state[2]), .I2(state[0]), 
            .I3(n3_adj_1353), .O(state_3__N_1123[0]));
    defparam i3861_3_lut_4_lut.LUT_INIT = 16'h1f0e;
    SB_CARRY counter_1437_add_4_8 (.CI(n12183), .I0(VCC_net), .I1(counter[6]), 
            .CO(n12184));
    SB_LUT4 counter_1437_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[5]), 
            .I3(n12182), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1437_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1186_7 (.CI(n12141), .I0(multi_byte_counter[5]), .I1(n2484[4]), 
            .CO(n12142));
    SB_LUT4 add_1186_6_lut (.I0(GND_net), .I1(multi_byte_counter[4]), .I2(n2484[4]), 
            .I3(n12140), .O(n315[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1186_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1186_6 (.CI(n12140), .I0(multi_byte_counter[4]), .I1(n2484[4]), 
            .CO(n12141));
    SB_CARRY counter_1437_add_4_7 (.CI(n12182), .I0(VCC_net), .I1(counter[5]), 
            .CO(n12183));
    SB_LUT4 add_1186_5_lut (.I0(GND_net), .I1(multi_byte_counter[3]), .I2(n2484[4]), 
            .I3(n12139), .O(n315[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1186_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1437_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[4]), 
            .I3(n12181), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1437_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1437_add_4_6 (.CI(n12181), .I0(VCC_net), .I1(counter[4]), 
            .CO(n12182));
    SB_CARRY add_1186_5 (.CI(n12139), .I0(multi_byte_counter[3]), .I1(n2484[4]), 
            .CO(n12140));
    SB_LUT4 counter_1437_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[3]), 
            .I3(n12180), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1437_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1437_add_4_5 (.CI(n12180), .I0(VCC_net), .I1(counter[3]), 
            .CO(n12181));
    SB_LUT4 counter_1437_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[2]), 
            .I3(n12179), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1437_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1186_4_lut (.I0(GND_net), .I1(multi_byte_counter[2]), .I2(n2484[4]), 
            .I3(n12138), .O(n315[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1186_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1437_add_4_4 (.CI(n12179), .I0(VCC_net), .I1(counter[2]), 
            .CO(n12180));
    SB_CARRY add_1186_4 (.CI(n12138), .I0(multi_byte_counter[2]), .I1(n2484[4]), 
            .CO(n12139));
    SB_LUT4 counter_1437_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[1]), 
            .I3(n12178), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1437_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1437_add_4_3 (.CI(n12178), .I0(VCC_net), .I1(counter[1]), 
            .CO(n12179));
    SB_LUT4 add_1186_3_lut (.I0(GND_net), .I1(multi_byte_counter[1]), .I2(n2484[4]), 
            .I3(n12137), .O(n315[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1186_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1437_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1437_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1186_3 (.CI(n12137), .I0(multi_byte_counter[1]), .I1(n2484[4]), 
            .CO(n12138));
    SB_LUT4 add_1186_2_lut (.I0(GND_net), .I1(multi_byte_counter[0]), .I2(n2484[4]), 
            .I3(GND_net), .O(n315[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1186_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1186_2 (.CI(GND_net), .I0(multi_byte_counter[0]), .I1(n2484[4]), 
            .CO(n12137));
    SB_CARRY counter_1437_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n12178));
    SB_LUT4 mux_1164_i16_3_lut (.I0(tx_addr_byte[7]), .I1(tx_shift_reg[14]), 
            .I2(n2407), .I3(GND_net), .O(n2408[15]));   // src/spi.v(88[9] 219[16])
    defparam mux_1164_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE tx_shift_reg_i0_i7 (.Q(tx_shift_reg[7]), .C(SLM_CLK_c), .E(n4837), 
            .D(n2408[7]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i8 (.Q(tx_shift_reg[8]), .C(SLM_CLK_c), .E(n4837), 
            .D(n2408[8]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i9 (.Q(tx_shift_reg[9]), .C(SLM_CLK_c), .E(n4837), 
            .D(n2408[9]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i10 (.Q(tx_shift_reg[10]), .C(SLM_CLK_c), .E(n4837), 
            .D(n2408[10]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i11 (.Q(tx_shift_reg[11]), .C(SLM_CLK_c), .E(n4837), 
            .D(n2408[11]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i12 (.Q(tx_shift_reg[12]), .C(SLM_CLK_c), .E(n4837), 
            .D(n2408[12]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i13 (.Q(tx_shift_reg[13]), .C(SLM_CLK_c), .E(n4837), 
            .D(n2408[13]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i14 (.Q(tx_shift_reg[14]), .C(SLM_CLK_c), .E(n4837), 
            .D(n2408[14]));   // src/spi.v(76[8] 221[4])
    SB_DFFESR counter_1437__i0 (.Q(counter[0]), .C(SLM_CLK_c), .E(n4912), 
            .D(n45[0]), .R(n5394));   // src/spi.v(183[28:41])
    SB_DFFESR multi_byte_counter_i0 (.Q(multi_byte_counter[0]), .C(SLM_CLK_c), 
            .E(n5054), .D(n315[0]), .R(n5383));   // src/spi.v(76[8] 221[4])
    SB_DFFESR counter_1437__i9 (.Q(counter[9]), .C(SLM_CLK_c), .E(n4912), 
            .D(n45[9]), .R(n5394));   // src/spi.v(183[28:41])
    SB_LUT4 mux_1164_i3_3_lut (.I0(\tx_data_byte[2] ), .I1(tx_shift_reg[1]), 
            .I2(n2407), .I3(GND_net), .O(n2408[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_1164_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS counter_1437__i8 (.Q(counter[8]), .C(SLM_CLK_c), .E(n4912), 
            .D(n45[8]), .S(n5394));   // src/spi.v(183[28:41])
    SB_LUT4 mux_1164_i4_3_lut (.I0(\tx_data_byte[3] ), .I1(tx_shift_reg[2]), 
            .I2(n2407), .I3(GND_net), .O(n2408[3]));   // src/spi.v(88[9] 219[16])
    defparam mux_1164_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR counter_1437__i7 (.Q(counter[7]), .C(SLM_CLK_c), .E(n4912), 
            .D(n45[7]), .R(n5394));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1437__i6 (.Q(counter[6]), .C(SLM_CLK_c), .E(n4912), 
            .D(n45[6]), .R(n5394));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1437__i5 (.Q(counter[5]), .C(SLM_CLK_c), .E(n4912), 
            .D(n45[5]), .R(n5394));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1437__i4 (.Q(counter[4]), .C(SLM_CLK_c), .E(n4912), 
            .D(n45[4]), .R(n5394));   // src/spi.v(183[28:41])
    SB_LUT4 mux_1164_i5_3_lut (.I0(\tx_data_byte[4] ), .I1(tx_shift_reg[3]), 
            .I2(n2407), .I3(GND_net), .O(n2408[4]));   // src/spi.v(88[9] 219[16])
    defparam mux_1164_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE state_i1 (.Q(state[1]), .C(SLM_CLK_c), .E(n12890), .D(state_3__N_1123[1]));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i2 (.Q(state[2]), .C(SLM_CLK_c), .E(n12889), .D(state_3__N_1123[2]));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i3 (.Q(state[3]), .C(SLM_CLK_c), .E(n19_adj_1354), .D(state_3__N_1123[3]));   // src/spi.v(76[8] 221[4])
    SB_DFF byte_recv_92_i3 (.Q(spi_rx_byte_ready), .C(SLM_CLK_c), .D(n1140[2]));   // src/spi.v(88[9] 219[16])
    SB_DFF byte_recv_92_i1 (.Q(SCK_c_0), .C(SLM_CLK_c), .D(n1140[0]));   // src/spi.v(88[9] 219[16])
    SB_LUT4 i10891_2_lut (.I0(state[0]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n13000));
    defparam i10891_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut (.I0(state[3]), .I1(n19), .I2(state[1]), .I3(GND_net), 
            .O(n12820));
    defparam i2_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i10895_2_lut (.I0(state[1]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n13004));
    defparam i10895_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(n13004), .I1(state[3]), .I2(spi_start_transfer_r), 
            .I3(state[0]), .O(n4896));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(state[3]), .I1(n4896), .I2(n19), .I3(state[0]), 
            .O(n6));
    defparam i2_4_lut.LUT_INIT = 16'hcc4c;
    SB_LUT4 i3_4_lut (.I0(n13004), .I1(n6), .I2(n5062), .I3(state[3]), 
            .O(n16230));
    defparam i3_4_lut.LUT_INIT = 16'h40c0;
    SB_LUT4 i12337_3_lut (.I0(counter[4]), .I1(n12829), .I2(n4570), .I3(GND_net), 
            .O(n4884));   // src/spi.v(88[9] 219[16])
    defparam i12337_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i2_3_lut_adj_37 (.I0(counter[1]), .I1(counter[3]), .I2(counter[2]), 
            .I3(GND_net), .O(n4705));   // src/spi.v(141[21:41])
    defparam i2_3_lut_adj_37.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_2_lut (.I0(multi_byte_counter[2]), .I1(multi_byte_counter[4]), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // src/spi.v(208[21:52])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(multi_byte_counter[3]), .I1(multi_byte_counter[1]), 
            .I2(multi_byte_counter[5]), .I3(multi_byte_counter[7]), .O(n14_adj_1355));   // src/spi.v(208[21:52])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(multi_byte_counter[0]), .I1(n14_adj_1355), .I2(n10), 
            .I3(multi_byte_counter[6]), .O(n2484[4]));   // src/spi.v(208[21:52])
    defparam i7_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i2_2_lut_adj_38 (.I0(counter[7]), .I1(counter[5]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_1356));   // src/spi.v(141[21:41])
    defparam i2_2_lut_adj_38.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_39 (.I0(counter[4]), .I1(counter[6]), .I2(counter[8]), 
            .I3(counter[9]), .O(n14_adj_1357));   // src/spi.v(141[21:41])
    defparam i6_4_lut_adj_39.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_40 (.I0(counter[0]), .I1(n14_adj_1357), .I2(n10_adj_1356), 
            .I3(n4705), .O(n19));   // src/spi.v(141[21:41])
    defparam i7_4_lut_adj_40.LUT_INIT = 16'hfffd;
    SB_LUT4 i12270_3_lut (.I0(n2484[4]), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n14298));   // src/spi.v(88[9] 219[16])
    defparam i12270_3_lut.LUT_INIT = 16'hc4c4;
    SB_LUT4 mux_380_Mux_1_i7_4_lut (.I0(state[0]), .I1(state[2]), .I2(n19), 
            .I3(state[1]), .O(n7));   // src/spi.v(88[9] 219[16])
    defparam mux_380_Mux_1_i7_4_lut.LUT_INIT = 16'h02dd;
    SB_LUT4 mux_380_Mux_1_i15_4_lut (.I0(n7), .I1(n14298), .I2(state[3]), 
            .I3(state[2]), .O(n1140[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_380_Mux_1_i15_4_lut.LUT_INIT = 16'hfaca;
    SB_DFFESR counter_1437__i3 (.Q(counter[3]), .C(SLM_CLK_c), .E(n4912), 
            .D(n45[3]), .R(n5394));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1437__i2 (.Q(counter[2]), .C(SLM_CLK_c), .E(n4912), 
            .D(n45[2]), .R(n5394));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1437__i1 (.Q(counter[1]), .C(SLM_CLK_c), .E(n4912), 
            .D(n45[1]), .R(n5394));   // src/spi.v(183[28:41])
    SB_DFF Rx_Recv_Byte_i0 (.Q(rx_buf_byte[0]), .C(SLM_CLK_c), .D(n5578));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i12216_2_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(state[2]), 
            .I3(GND_net), .O(n14305));
    defparam i12216_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(state[2]), 
            .I3(GND_net), .O(n24));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 mux_1164_i6_3_lut (.I0(\tx_data_byte[5] ), .I1(tx_shift_reg[4]), 
            .I2(n2407), .I3(GND_net), .O(n2408[5]));   // src/spi.v(88[9] 219[16])
    defparam mux_1164_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_41 (.I0(counter[0]), .I1(counter[1]), .I2(counter[2]), 
            .I3(counter[3]), .O(n12829));
    defparam i3_4_lut_adj_41.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_42 (.I0(state[3]), .I1(state[1]), .I2(state[0]), 
            .I3(state[2]), .O(n4));
    defparam i1_4_lut_adj_42.LUT_INIT = 16'h4046;
    SB_LUT4 i1_3_lut_adj_43 (.I0(counter[4]), .I1(n4), .I2(n12829), .I3(GND_net), 
            .O(n2407));
    defparam i1_3_lut_adj_43.LUT_INIT = 16'h4040;
    SB_LUT4 i1_4_lut_adj_44 (.I0(n12829), .I1(state[3]), .I2(counter[4]), 
            .I3(state[1]), .O(n16));   // src/spi.v(88[9] 219[16])
    defparam i1_4_lut_adj_44.LUT_INIT = 16'hf5c4;
    SB_LUT4 i30_4_lut (.I0(spi_start_transfer_r), .I1(state[3]), .I2(state[1]), 
            .I3(state[0]), .O(n24_adj_1358));   // src/spi.v(88[9] 219[16])
    defparam i30_4_lut.LUT_INIT = 16'hcfc1;
    SB_LUT4 mux_1164_i7_3_lut (.I0(\tx_data_byte[6] ), .I1(tx_shift_reg[5]), 
            .I2(n2407), .I3(GND_net), .O(n2408[6]));   // src/spi.v(88[9] 219[16])
    defparam mux_1164_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(counter[0]), .I1(counter[1]), .I2(counter[3]), 
            .I3(counter[2]), .O(n8));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12219_2_lut_4_lut (.I0(state[2]), .I1(state[0]), .I2(state[1]), 
            .I3(n8), .O(n14272));   // src/spi.v(88[9] 219[16])
    defparam i12219_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 mux_380_Mux_2_i15_4_lut_4_lut (.I0(state[0]), .I1(state[2]), 
            .I2(state[3]), .I3(state[1]), .O(n1140[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_380_Mux_2_i15_4_lut_4_lut.LUT_INIT = 16'h1008;
    SB_LUT4 i10927_3_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(spi_start_transfer_r), 
            .I3(state[2]), .O(n13036));
    defparam i10927_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12378_3_lut_4_lut (.I0(state[2]), .I1(state[0]), .I2(n24_adj_1358), 
            .I3(n16), .O(n4837));   // src/spi.v(88[9] 219[16])
    defparam i12378_3_lut_4_lut.LUT_INIT = 16'h000d;
    SB_LUT4 i3099_4_lut_4_lut (.I0(state[2]), .I1(state[0]), .I2(state[1]), 
            .I3(state[3]), .O(n4570));   // src/spi.v(88[9] 219[16])
    defparam i3099_4_lut_4_lut.LUT_INIT = 16'hfe2f;
    SB_LUT4 mux_56_Mux_1_i15_3_lut_4_lut (.I0(state[0]), .I1(state[1]), 
            .I2(state[3]), .I3(n7_adj_1359), .O(state_3__N_1123[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_1_i15_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i2_2_lut_4_lut (.I0(state[3]), .I1(n19), .I2(state[1]), .I3(n13000), 
            .O(n5062));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 mux_56_Mux_1_i7_4_lut (.I0(n3), .I1(n14309), .I2(state[2]), 
            .I3(state[1]), .O(n7_adj_1359));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_1_i7_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i12275_2_lut (.I0(n19), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n14309));   // src/spi.v(88[9] 219[16])
    defparam i12275_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_3_lut_adj_45 (.I0(state[3]), .I1(n12888), .I2(n24), .I3(GND_net), 
            .O(n12890));
    defparam i1_3_lut_adj_45.LUT_INIT = 16'h4c4c;
    SB_LUT4 i1_3_lut_adj_46 (.I0(n4896), .I1(state[2]), .I2(n12820), .I3(GND_net), 
            .O(n12888));
    defparam i1_3_lut_adj_46.LUT_INIT = 16'ha8a8;
    SB_LUT4 mux_56_Mux_2_i15_4_lut (.I0(n3_adj_1360), .I1(state[2]), .I2(state[3]), 
            .I3(state[0]), .O(state_3__N_1123[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_2_i15_4_lut.LUT_INIT = 16'hc2ce;
    SB_LUT4 mux_56_Mux_2_i3_3_lut (.I0(multi_byte_spi_trans_flag_r), .I1(state[0]), 
            .I2(state[1]), .I3(GND_net), .O(n3_adj_1360));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_2_i3_3_lut.LUT_INIT = 16'hc2c2;
    SB_LUT4 i1_2_lut (.I0(n5062), .I1(n12888), .I2(GND_net), .I3(GND_net), 
            .O(n12889));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_56_Mux_3_i15_4_lut (.I0(n14305), .I1(state[1]), .I2(state[3]), 
            .I3(n2484[4]), .O(state_3__N_1123[3]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_3_i15_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i12315_4_lut (.I0(n22), .I1(n13036), .I2(n24), .I3(state[3]), 
            .O(n19_adj_1354));
    defparam i12315_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i1_2_lut_adj_47 (.I0(n19), .I1(n21), .I2(GND_net), .I3(GND_net), 
            .O(n22));
    defparam i1_2_lut_adj_47.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_48 (.I0(counter[4]), .I1(n14271), .I2(n14272), 
            .I3(state[3]), .O(n1140[0]));   // src/spi.v(88[9] 219[16])
    defparam i1_4_lut_adj_48.LUT_INIT = 16'ha088;
    SB_LUT4 i12276_4_lut (.I0(n8), .I1(state[1]), .I2(state[0]), .I3(state[2]), 
            .O(n14271));   // src/spi.v(88[9] 219[16])
    defparam i12276_4_lut.LUT_INIT = 16'hc08c;
    SB_LUT4 i12225_2_lut_3_lut (.I0(n19), .I1(state[0]), .I2(state[2]), 
            .I3(GND_net), .O(n14300));
    defparam i12225_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i2500_4_lut_4_lut (.I0(state[2]), .I1(state[3]), .I2(state[0]), 
            .I3(state[1]), .O(n3963));   // src/spi.v(88[9] 219[16])
    defparam i2500_4_lut_4_lut.LUT_INIT = 16'hffbd;
    SB_LUT4 i1_3_lut_4_lut (.I0(n2484[4]), .I1(state[0]), .I2(state[2]), 
            .I3(state[1]), .O(n4776));   // src/spi.v(88[9] 219[16])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfdfc;
>>>>>>> Stashed changes
>>>>>>> master
    
endmodule

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Mar 10 2020 15:49:36

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    SOUT : in std_logic;
    SCK : out std_logic;
    FIFO_D31 : in std_logic;
    FIFO_D20 : in std_logic;
    FIFO_D13 : in std_logic;
    FIFO_D1 : in std_logic;
    FIFO_CLK : in std_logic;
    FIFO_BE2 : in std_logic;
    DATA15 : out std_logic;
    DATA4 : out std_logic;
    DATA23 : out std_logic;
    RST : out std_logic;
    FIFO_D4 : in std_logic;
    FIFO_D14 : in std_logic;
    UART_TX : out std_logic;
    DATA10 : out std_logic;
    DATA28 : out std_logic;
    DATA19 : out std_logic;
    SDAT : out std_logic;
    FT_SIWU : out std_logic;
    DATA0 : out std_logic;
    FT_WR : out std_logic;
    FIFO_D27 : in std_logic;
    FIFO_D10 : in std_logic;
    FIFO_D0 : in std_logic;
    FIFO_BE3 : in std_logic;
    DEBUG_0 : out std_logic;
    FIFO_D9 : in std_logic;
    DATA14 : out std_logic;
    UPDATE : out std_logic;
    RESET : out std_logic;
    FIFO_D21 : in std_logic;
    FIFO_D12 : in std_logic;
    FIFO_BE1 : in std_logic;
    DEBUG_6 : out std_logic;
    DATA5 : out std_logic;
    DATA24 : out std_logic;
    SEN : out std_logic;
    FIFO_D7 : in std_logic;
    FIFO_D15 : in std_logic;
    ICE_CREST : out std_logic;
    FIFO_D23 : in std_logic;
    DATA3 : out std_logic;
    DATA22 : out std_logic;
    DATA13 : out std_logic;
    INVERT : out std_logic;
    FT_RD : out std_logic;
    FIFO_D5 : in std_logic;
    FIFO_D24 : in std_logic;
    FIFO_D17 : in std_logic;
    DSR : out std_logic;
    DEBUG_3 : out std_logic;
    DATA29 : out std_logic;
    DATA18 : out std_logic;
    ICE_SYSCLK : in std_logic;
    ICE_CLK : out std_logic;
    DATA20 : out std_logic;
    DATA11 : out std_logic;
    DATA1 : out std_logic;
    VALID : out std_logic;
    SYNC : out std_logic;
    FIFO_D3 : in std_logic;
    FIFO_D26 : in std_logic;
    FIFO_D11 : in std_logic;
    DEBUG_1 : out std_logic;
    DATA8 : out std_logic;
    DATA31 : out std_logic;
    DATA27 : out std_logic;
    CTS : out std_logic;
    FIFO_D8 : in std_logic;
    FIFO_D18 : in std_logic;
    DEBUG_8 : out std_logic;
    DCD : out std_logic;
    DATA17 : out std_logic;
    SLM_CLK : out std_logic;
    DATA6 : out std_logic;
    DATA25 : out std_logic;
    ICE_CDONE : out std_logic;
    FIFO_D6 : in std_logic;
    FIFO_D29 : in std_logic;
    UART_RX : in std_logic;
    FIFO_D22 : in std_logic;
    FIFO_BE0 : in std_logic;
    DEBUG_5 : out std_logic;
    DATA12 : out std_logic;
    DTR : out std_logic;
    DATA21 : out std_logic;
    DATA2 : out std_logic;
    FIFO_D25 : in std_logic;
    FIFO_D2 : in std_logic;
    FIFO_D16 : in std_logic;
    DEBUG_2 : out std_logic;
    DATA9 : out std_logic;
    DATA30 : out std_logic;
    FT_TXE : in std_logic;
    FR_RXF : in std_logic;
    FIFO_D19 : in std_logic;
    DEBUG_9 : out std_logic;
    DATA16 : out std_logic;
    FT_OE : out std_logic;
    DATA7 : out std_logic;
    DATA26 : out std_logic;
    FIFO_D30 : in std_logic;
    FIFO_D28 : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__20524\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17196\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17034\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16731\ : std_logic;
signal \N__16728\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16651\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16641\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16416\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14970\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14910\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14679\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14193\ : std_logic;
signal \N__14190\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13462\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13435\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \FT_RD_c\ : std_logic;
signal \FIFO_D19_c_19\ : std_logic;
signal \DATA19_c_19\ : std_logic;
signal \FIFO_D14_c_14\ : std_logic;
signal \DATA14_c_14\ : std_logic;
signal \FIFO_D30_c_30\ : std_logic;
signal \DATA30_c_30\ : std_logic;
signal \FIFO_D31_c_31\ : std_logic;
signal \DATA31_c_31\ : std_logic;
signal \FIFO_D11_c_11\ : std_logic;
signal \DATA11_c_11\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_0\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_0\ : std_logic;
signal rx_shift_reg_8 : std_logic;
signal rx_shift_reg_7 : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_3\ : std_logic;
signal \SOUT_c\ : std_logic;
signal rx_shift_reg_0 : std_logic;
signal \FIFO_D28_c_28\ : std_logic;
signal \DATA28_c_28\ : std_logic;
signal \SCK_c\ : std_logic;
signal \FIFO_D23_c_23\ : std_logic;
signal \DATA23_c_23\ : std_logic;
signal rx_buf_byte_0 : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_0\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n5666\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_0\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_2\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_3\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_5\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_5\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_3\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_3\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n5690\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_6\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_6\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n5696_cascade_\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_6\ : std_logic;
signal \mem_LUT_data_raw_r_6\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n5702\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_5\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_5\ : std_logic;
signal rx_shift_reg_6 : std_logic;
signal rx_buf_byte_5 : std_logic;
signal rx_shift_reg_4 : std_logic;
signal rx_buf_byte_3 : std_logic;
signal rx_shift_reg_1 : std_logic;
signal rx_shift_reg_2 : std_logic;
signal rx_shift_reg_3 : std_logic;
signal \SEN_c\ : std_logic;
signal \FIFO_D25_c_25\ : std_logic;
signal \DATA25_c_25\ : std_logic;
signal \FIFO_D29_c_29\ : std_logic;
signal \DATA29_c_29\ : std_logic;
signal rx_buf_byte_2 : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_2\ : std_logic;
signal fifo_temp_output_6 : std_logic;
signal \pc_tx.n3763_cascade_\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_2\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n5660\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_2\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_1\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_1\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_1\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n5672_cascade_\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n5678_cascade_\ : std_logic;
signal \mem_LUT_data_raw_r_4\ : std_logic;
signal \spi0.n480\ : std_logic;
signal \spi0.state_next_1_cascade_\ : std_logic;
signal \spi0.n481\ : std_logic;
signal \spi0.n482\ : std_logic;
signal \spi0.n483\ : std_logic;
signal \spi0.n484\ : std_logic;
signal \spi0.n485\ : std_logic;
signal \spi0.n490\ : std_logic;
signal \spi0.n488\ : std_logic;
signal \spi0.n487\ : std_logic;
signal \spi0.n486\ : std_logic;
signal rx_buf_byte_6 : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_6\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_7\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_7\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_4\ : std_logic;
signal \spi0.n14_cascade_\ : std_logic;
signal rx_shift_reg_5 : std_logic;
signal \rx_shift_reg_15__N_461\ : std_logic;
signal \spi0.n10\ : std_logic;
signal \spi0.spi_clk_counter_0\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \spi0.spi_clk_counter_1\ : std_logic;
signal \spi0.n4874\ : std_logic;
signal \spi0.spi_clk_counter_2\ : std_logic;
signal \spi0.n4875\ : std_logic;
signal \spi0.spi_clk_counter_3\ : std_logic;
signal \spi0.n4876\ : std_logic;
signal \spi0.spi_clk_counter_4\ : std_logic;
signal \spi0.n4877\ : std_logic;
signal \spi0.spi_clk_counter_5\ : std_logic;
signal \spi0.n4878\ : std_logic;
signal \spi0.spi_clk_counter_6\ : std_logic;
signal \spi0.n4879\ : std_logic;
signal \spi0.n4880\ : std_logic;
signal \spi0.spi_clk_counter_7\ : std_logic;
signal \FIFO_D18_c_18\ : std_logic;
signal \DATA18_c_18\ : std_logic;
signal \mem_LUT_data_raw_r_2\ : std_logic;
signal fifo_temp_output_4 : std_logic;
signal fifo_temp_output_2 : std_logic;
signal \r_Tx_Data_3\ : std_logic;
signal \r_Tx_Data_2\ : std_logic;
signal \r_Tx_Data_5\ : std_logic;
signal \r_Tx_Data_4\ : std_logic;
signal n5414 : std_logic;
signal \r_Tx_Data_6\ : std_logic;
signal \pc_tx.r_Bit_Index_1\ : std_logic;
signal \pc_tx.n5512_cascade_\ : std_logic;
signal \pc_tx.n5511\ : std_logic;
signal \pc_tx.r_Bit_Index_2\ : std_logic;
signal \pc_tx.n5654_cascade_\ : std_logic;
signal \pc_tx.n5509\ : std_logic;
signal \pc_tx.o_Tx_Serial_N_354_cascade_\ : std_logic;
signal \pc_tx.n3_adj_632\ : std_logic;
signal \pc_tx.n5486\ : std_logic;
signal \n2366_cascade_\ : std_logic;
signal \r_Tx_Data_7\ : std_logic;
signal \pc_tx.r_Bit_Index_0\ : std_logic;
signal \pc_tx.n5508\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_4\ : std_logic;
signal \mem_LUT_data_raw_r_3\ : std_logic;
signal fifo_temp_output_3 : std_logic;
signal \mem_LUT_data_raw_r_0\ : std_logic;
signal rx_buf_byte_1 : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_1\ : std_logic;
signal \r_Tx_Data_1\ : std_logic;
signal fifo_temp_output_0 : std_logic;
signal n2366 : std_logic;
signal \r_Tx_Data_0\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_4\ : std_logic;
signal \spi0.n2120_cascade_\ : std_logic;
signal \spi0.n5552\ : std_logic;
signal \spi0.n5552_cascade_\ : std_logic;
signal \spi0.state_next_2_cascade_\ : std_logic;
signal \spi0.n4_cascade_\ : std_logic;
signal \spi0.n492\ : std_logic;
signal \spi0.n491\ : std_logic;
signal \state_next_2__N_454\ : std_logic;
signal \spi0.n1005\ : std_logic;
signal \n982_cascade_\ : std_logic;
signal \spi0.state_next_1\ : std_logic;
signal \spi0.n495\ : std_logic;
signal \spi0.n4\ : std_logic;
signal \spi0.state_next_2__N_453\ : std_logic;
signal \spi0.state_next_2__N_452\ : std_logic;
signal \spi0.n5561_cascade_\ : std_logic;
signal \spi0.n25\ : std_logic;
signal \spi0.n13\ : std_logic;
signal n982 : std_logic;
signal \spi0.n2120\ : std_logic;
signal \spi0.n13_cascade_\ : std_logic;
signal \spi0.state_next_0\ : std_logic;
signal \mem_LUT_data_raw_r_5\ : std_logic;
signal fifo_temp_output_5 : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_7\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n5684\ : std_logic;
signal \mem_LUT_data_raw_r_1\ : std_logic;
signal fifo_temp_output_1 : std_logic;
signal \FIFO_D8_c_8\ : std_logic;
signal \DATA8_c_8\ : std_logic;
signal \spi0.CS_w\ : std_logic;
signal \spi0.n2715\ : std_logic;
signal \pc_tx.n5_cascade_\ : std_logic;
signal \pc_tx.n4905_cascade_\ : std_logic;
signal \pc_tx.r_SM_Main_2_N_322_1_cascade_\ : std_logic;
signal \pc_tx.n3763\ : std_logic;
signal \pc_tx.n2069\ : std_logic;
signal \pc_tx.n5484\ : std_logic;
signal \pc_tx.n6\ : std_logic;
signal \spi0.spi_clk\ : std_logic;
signal \n2446_cascade_\ : std_logic;
signal tx_shift_reg_4 : std_logic;
signal tx_shift_reg_8 : std_logic;
signal tx_shift_reg_3 : std_logic;
signal tx_shift_reg_9 : std_logic;
signal tx_shift_reg_10 : std_logic;
signal \INVspi0.tx_shift_reg_i8C_net\ : std_logic;
signal tx_shift_reg_5 : std_logic;
signal \n5462_cascade_\ : std_logic;
signal tx_shift_reg_6 : std_logic;
signal tx_shift_reg_7 : std_logic;
signal \INVspi0.tx_shift_reg_i6C_net\ : std_logic;
signal rx_buf_byte_7 : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_7\ : std_logic;
signal \r_SM_Main_2_N_325_0\ : std_logic;
signal rx_buf_byte_4 : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_4\ : std_logic;
signal \reset_all_w_N_61\ : std_logic;
signal reset_clk_counter_0 : std_logic;
signal \reset_all_w_N_61_cascade_\ : std_logic;
signal reset_clk_counter_1 : std_logic;
signal \n2_adj_670_cascade_\ : std_logic;
signal reset_clk_counter_2 : std_logic;
signal reset_clk_counter_3 : std_logic;
signal \FIFO_D26_c_26\ : std_logic;
signal \DATA26_c_26\ : std_logic;
signal \FIFO_D15_c_15\ : std_logic;
signal \DATA15_c_15\ : std_logic;
signal spi_busy : std_logic;
signal spi_busy_prev : std_logic;
signal \tx_fifo.lscc_fifo_inst.n4\ : std_logic;
signal spi_busy_falling_edge : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3\ : std_logic;
signal \pc_tx.r_Clock_Count_0\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \pc_tx.r_Clock_Count_1\ : std_logic;
signal \pc_tx.n4865\ : std_logic;
signal \pc_tx.r_Clock_Count_2\ : std_logic;
signal \pc_tx.n4866\ : std_logic;
signal \pc_tx.r_Clock_Count_3\ : std_logic;
signal \pc_tx.n4867\ : std_logic;
signal \pc_tx.r_Clock_Count_4\ : std_logic;
signal \pc_tx.n4868\ : std_logic;
signal \pc_tx.r_Clock_Count_5\ : std_logic;
signal \pc_tx.n4869\ : std_logic;
signal \pc_tx.r_Clock_Count_6\ : std_logic;
signal \pc_tx.n4870\ : std_logic;
signal \pc_tx.r_Clock_Count_7\ : std_logic;
signal \pc_tx.n4871\ : std_logic;
signal \pc_tx.n4872\ : std_logic;
signal \pc_tx.r_Clock_Count_8\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \pc_tx.n4873\ : std_logic;
signal \pc_tx.r_Clock_Count_9\ : std_logic;
signal \pc_tx.n2739\ : std_logic;
signal \DEBUG_9_c\ : std_logic;
signal tx_shift_reg_11 : std_logic;
signal tx_shift_reg_2 : std_logic;
signal tx_shift_reg_12 : std_logic;
signal tx_shift_reg_13 : std_logic;
signal tx_shift_reg_14 : std_logic;
signal n5462 : std_logic;
signal n2446 : std_logic;
signal tx_shift_reg_1 : std_logic;
signal \INVspi0.tx_shift_reg_i15C_net\ : std_logic;
signal tx_uart_active_flag : std_logic;
signal \n5454_cascade_\ : std_logic;
signal \RESET_c\ : std_logic;
signal \n15_adj_673_cascade_\ : std_logic;
signal n4892 : std_logic;
signal \tx_fifo.lscc_fifo_inst.rd_addr_r_2\ : std_logic;
signal n1 : std_logic;
signal \tx_fifo.lscc_fifo_inst.rd_fifo_en_w\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.rd_fifo_en_w_cascade_\ : std_logic;
signal \mem_LUT_data_raw_r_7\ : std_logic;
signal fifo_temp_output_7 : std_logic;
signal is_tx_fifo_full_flag : std_logic;
signal \FIFO_D27_c_27\ : std_logic;
signal \DATA27_c_27\ : std_logic;
signal \FIFO_D20_c_20\ : std_logic;
signal \DATA20_c_20\ : std_logic;
signal \FIFO_D13_c_13\ : std_logic;
signal \DATA13_c_13\ : std_logic;
signal tx_addr_byte_4 : std_logic;
signal \pc_rx.n5450\ : std_logic;
signal \pc_rx.n1\ : std_logic;
signal tx_addr_byte_1 : std_logic;
signal tx_addr_byte_5 : std_logic;
signal pc_data_rx_1 : std_logic;
signal tx_data_byte_1 : std_logic;
signal \pc_rx.n5452_cascade_\ : std_logic;
signal \pc_rx.n5478_cascade_\ : std_logic;
signal \pc_rx.n6\ : std_logic;
signal \pc_rx.n5488_cascade_\ : std_logic;
signal \pc_rx.r_SM_Main_2_N_252_0\ : std_logic;
signal \pc_rx.r_SM_Main_2_N_252_0_cascade_\ : std_logic;
signal \pc_rx.n6_adj_635\ : std_logic;
signal tx_data_byte_7 : std_logic;
signal tx_addr_byte_7 : std_logic;
signal state_reg_0 : std_logic;
signal tx_addr_byte_2 : std_logic;
signal wr_addr_p1_w_2 : std_logic;
signal \wr_addr_p1_w_2_cascade_\ : std_logic;
signal wr_fifo_en_w : std_logic;
signal \tx_fifo.lscc_fifo_inst.n2\ : std_logic;
signal rd_addr_r_1 : std_logic;
signal \n32_cascade_\ : std_logic;
signal fifo_write_cmd : std_logic;
signal wr_addr_r_2 : std_logic;
signal rd_addr_p1_w_1 : std_logic;
signal rd_addr_p1_w_2 : std_logic;
signal wr_addr_r_1 : std_logic;
signal \n5474_cascade_\ : std_logic;
signal n24_adj_674 : std_logic;
signal wr_addr_r_0 : std_logic;
signal n4_adj_675 : std_logic;
signal n2545 : std_logic;
signal \tx_fifo.lscc_fifo_inst.rd_fifo_en_prev_r\ : std_logic;
signal \FIFO_D24_c_24\ : std_logic;
signal \DATA24_c_24\ : std_logic;
signal \FIFO_D5_c_5\ : std_logic;
signal \DATA5_c_5\ : std_logic;
signal \FIFO_D6_c_6\ : std_logic;
signal \DATA6_c_6\ : std_logic;
signal n4 : std_logic;
signal tx_data_byte_4 : std_logic;
signal \n2468_cascade_\ : std_logic;
signal pc_data_rx_5 : std_logic;
signal tx_data_byte_5 : std_logic;
signal n2468 : std_logic;
signal pc_data_rx_4 : std_logic;
signal \pc_rx.n3803\ : std_logic;
signal \n2475_cascade_\ : std_logic;
signal pc_data_rx_7 : std_logic;
signal n2475 : std_logic;
signal pc_data_rx_3 : std_logic;
signal \pc_rx.n2465_cascade_\ : std_logic;
signal \pc_rx.n4887_cascade_\ : std_logic;
signal \r_SM_Main_2_N_246_2_cascade_\ : std_logic;
signal \pc_rx.n2429\ : std_logic;
signal \pc_rx.n2429_cascade_\ : std_logic;
signal \bfn_13_6_0_\ : std_logic;
signal \pc_rx.n4807\ : std_logic;
signal \pc_rx.r_Clock_Count_2\ : std_logic;
signal \pc_rx.n4808\ : std_logic;
signal \pc_rx.r_Clock_Count_3\ : std_logic;
signal \pc_rx.n4809\ : std_logic;
signal \pc_rx.n4810\ : std_logic;
signal \pc_rx.r_Clock_Count_5\ : std_logic;
signal \pc_rx.n4811\ : std_logic;
signal \pc_rx.r_Clock_Count_6\ : std_logic;
signal \pc_rx.n4812\ : std_logic;
signal \pc_rx.r_Clock_Count_7\ : std_logic;
signal \pc_rx.n4813\ : std_logic;
signal \pc_rx.n4814\ : std_logic;
signal \pc_rx.r_Clock_Count_8\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \pc_rx.n4815\ : std_logic;
signal \pc_rx.r_Clock_Count_9\ : std_logic;
signal \pc_rx.n2566\ : std_logic;
signal \pc_rx.n2705\ : std_logic;
signal state_reg_2 : std_logic;
signal state_reg_1 : std_logic;
signal tx_shift_reg_0 : std_logic;
signal \INVspi0.tx_shift_reg_i0C_net\ : std_logic;
signal n989 : std_logic;
signal \bluejay_data_inst.n1040_cascade_\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_7_N_122_3_cascade_\ : std_logic;
signal \bluejay_data_inst.n8_adj_656_cascade_\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_7_N_122_3\ : std_logic;
signal \bluejay_data_inst.n1041_cascade_\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_7_N_122_2_cascade_\ : std_logic;
signal \bluejay_data_inst.n18_cascade_\ : std_logic;
signal \bluejay_data_inst.n20\ : std_logic;
signal \bluejay_data_inst.n1675\ : std_logic;
signal \FIFO_D1_c_1\ : std_logic;
signal \DATA1_c_1\ : std_logic;
signal \FIFO_D21_c_21\ : std_logic;
signal \DATA21_c_21\ : std_logic;
signal \pc_rx.n5522_cascade_\ : std_logic;
signal \n5482_cascade_\ : std_logic;
signal n3753 : std_logic;
signal \r_SM_Main_2_N_246_2\ : std_logic;
signal \r_SM_Main_0\ : std_logic;
signal \r_SM_Main_2\ : std_logic;
signal \n2502_cascade_\ : std_logic;
signal \r_SM_Main_1\ : std_logic;
signal \pc_rx.r_Clock_Count_1\ : std_logic;
signal \pc_rx.r_Clock_Count_4\ : std_logic;
signal \pc_rx.r_Clock_Count_0\ : std_logic;
signal \pc_rx.n4\ : std_logic;
signal pc_data_rx_0 : std_logic;
signal \usb_to_bluejay_if_inst.n5438_cascade_\ : std_logic;
signal tx_addr_byte_6 : std_logic;
signal tx_data_byte_6 : std_logic;
signal n3672 : std_logic;
signal pc_data_rx_6 : std_logic;
signal n4_adj_666 : std_logic;
signal n2471 : std_logic;
signal pc_data_rx_2 : std_logic;
signal tx_data_byte_2 : std_logic;
signal tx_data_byte_3 : std_logic;
signal tx_addr_byte_3 : std_logic;
signal tx_data_byte_0 : std_logic;
signal tx_addr_byte_0 : std_logic;
signal \bluejay_data_inst.n5531\ : std_logic;
signal \bluejay_data_inst.n19\ : std_logic;
signal fifo_read_cmd : std_logic;
signal is_fifo_empty_flag : std_logic;
signal rd_addr_r_0 : std_logic;
signal \FIFO_D10_c_10\ : std_logic;
signal \DATA10_c_10\ : std_logic;
signal \FIFO_D9_c_9\ : std_logic;
signal \DATA9_c_9\ : std_logic;
signal \FIFO_D16_c_16\ : std_logic;
signal \DATA16_c_16\ : std_logic;
signal \pc_rx.r_Bit_Index_2\ : std_logic;
signal \r_Bit_Index_0\ : std_logic;
signal \pc_rx.r_Bit_Index_1\ : std_logic;
signal n5482 : std_logic;
signal \pc_rx.n2676\ : std_logic;
signal debug_led3 : std_logic;
signal uart_rx_complete_prev : std_logic;
signal n5_adj_667 : std_logic;
signal start_transfer_edge : std_logic;
signal \usb_to_bluejay_if_inst.n5400_cascade_\ : std_logic;
signal \usb_to_bluejay_if_inst.n2527_cascade_\ : std_logic;
signal spi_start_transfer_r : std_logic;
signal start_transfer_prev : std_logic;
signal data_in_fifo_prev : std_logic;
signal \usb_to_bluejay_if_inst.n4136_cascade_\ : std_logic;
signal \usb_to_bluejay_if_inst.n2492_cascade_\ : std_logic;
signal \usb_to_bluejay_if_inst.n2492\ : std_logic;
signal \usb_to_bluejay_if_inst.n4963\ : std_logic;
signal \usb_to_bluejay_if_inst.n3\ : std_logic;
signal \usb_to_bluejay_if_inst.state_timeout_counter_7__N_178_cascade_\ : std_logic;
signal \usb_to_bluejay_if_inst.n5400\ : std_logic;
signal \usb_to_bluejay_if_inst.n2562_cascade_\ : std_logic;
signal \usb_to_bluejay_if_inst.n2564\ : std_logic;
signal \usb_to_bluejay_if_inst.n2564_cascade_\ : std_logic;
signal \usb_to_bluejay_if_inst.n2706\ : std_logic;
signal \bfn_15_8_0_\ : std_logic;
signal \bluejay_data_inst.v_counter_0\ : std_logic;
signal \bluejay_data_inst.n1476\ : std_logic;
signal \bluejay_data_inst.n1109\ : std_logic;
signal \bluejay_data_inst.n4847\ : std_logic;
signal \bluejay_data_inst.v_counter_1\ : std_logic;
signal \bluejay_data_inst.n1108\ : std_logic;
signal \bluejay_data_inst.n4848\ : std_logic;
signal \bluejay_data_inst.v_counter_2\ : std_logic;
signal \bluejay_data_inst.n1107\ : std_logic;
signal \bluejay_data_inst.n4849\ : std_logic;
signal \bluejay_data_inst.v_counter_3\ : std_logic;
signal \bluejay_data_inst.n1106\ : std_logic;
signal \bluejay_data_inst.n4850\ : std_logic;
signal \bluejay_data_inst.v_counter_4\ : std_logic;
signal \bluejay_data_inst.n1105\ : std_logic;
signal \bluejay_data_inst.n4851\ : std_logic;
signal \bluejay_data_inst.v_counter_5\ : std_logic;
signal \bluejay_data_inst.n1104\ : std_logic;
signal \bluejay_data_inst.n4852\ : std_logic;
signal \bluejay_data_inst.v_counter_6\ : std_logic;
signal \bluejay_data_inst.n1103\ : std_logic;
signal \bluejay_data_inst.n4853\ : std_logic;
signal \bluejay_data_inst.n4854\ : std_logic;
signal \bluejay_data_inst.v_counter_7\ : std_logic;
signal \bluejay_data_inst.n1102\ : std_logic;
signal \bfn_15_9_0_\ : std_logic;
signal \bluejay_data_inst.v_counter_8\ : std_logic;
signal \bluejay_data_inst.n1101\ : std_logic;
signal \bluejay_data_inst.n4855\ : std_logic;
signal \bluejay_data_inst.v_counter_9\ : std_logic;
signal \bluejay_data_inst.n1100\ : std_logic;
signal \bluejay_data_inst.n4856\ : std_logic;
signal \bluejay_data_inst.v_counter_10\ : std_logic;
signal \bluejay_data_inst.n4857\ : std_logic;
signal \bluejay_data_inst.n1099\ : std_logic;
signal \bluejay_data_inst.n1054_cascade_\ : std_logic;
signal \bluejay_data_inst.n1373\ : std_logic;
signal \n5_cascade_\ : std_logic;
signal \bluejay_data_inst.n5524\ : std_logic;
signal \bluejay_data_inst.n1432\ : std_logic;
signal \FIFO_D3_c_3\ : std_logic;
signal \DATA3_c_3\ : std_logic;
signal \n3_adj_669_cascade_\ : std_logic;
signal \FIFO_D12_c_12\ : std_logic;
signal \DATA12_c_12\ : std_logic;
signal uart_rx_complete_rising_edge : std_logic;
signal even_byte_flag : std_logic;
signal \bfn_16_5_0_\ : std_logic;
signal \usb_to_bluejay_if_inst.n4800\ : std_logic;
signal \usb_to_bluejay_if_inst.n4801\ : std_logic;
signal \usb_to_bluejay_if_inst.state_timeout_counter_3\ : std_logic;
signal \usb_to_bluejay_if_inst.n82\ : std_logic;
signal \usb_to_bluejay_if_inst.n4802\ : std_logic;
signal \usb_to_bluejay_if_inst.n4803\ : std_logic;
signal \usb_to_bluejay_if_inst.n81\ : std_logic;
signal \usb_to_bluejay_if_inst.state_timeout_counter_5\ : std_logic;
signal \usb_to_bluejay_if_inst.n83\ : std_logic;
signal \usb_to_bluejay_if_inst.n4804\ : std_logic;
signal \usb_to_bluejay_if_inst.state_timeout_counter_6\ : std_logic;
signal \usb_to_bluejay_if_inst.n4805\ : std_logic;
signal \usb_to_bluejay_if_inst.n4806\ : std_logic;
signal \usb_to_bluejay_if_inst.state_timeout_counter_7\ : std_logic;
signal \usb_to_bluejay_if_inst.n2527\ : std_logic;
signal \usb_to_bluejay_if_inst.n4120\ : std_logic;
signal \usb_to_bluejay_if_inst.state_timeout_counter_2\ : std_logic;
signal \usb_to_bluejay_if_inst.state_timeout_counter_1\ : std_logic;
signal \usb_to_bluejay_if_inst.state_timeout_counter_4\ : std_logic;
signal \usb_to_bluejay_if_inst.state_timeout_counter_0\ : std_logic;
signal \usb_to_bluejay_if_inst.n12_cascade_\ : std_logic;
signal \usb_to_bluejay_if_inst.n13\ : std_logic;
signal n11 : std_logic;
signal \n11_cascade_\ : std_logic;
signal state_2_adj_657 : std_logic;
signal state_1 : std_logic;
signal \usb_to_bluejay_if_inst.n82_adj_628_cascade_\ : std_logic;
signal \usb_to_bluejay_if_inst.state_timeout_counter_7__N_178\ : std_logic;
signal \usb_to_bluejay_if_inst.n2561\ : std_logic;
signal \pc_tx.r_SM_Main_0\ : std_logic;
signal \r_SM_Main_1_adj_660\ : std_logic;
signal \pc_tx.r_SM_Main_2_N_322_1\ : std_logic;
signal n10_adj_671 : std_logic;
signal n16_adj_672 : std_logic;
signal state_0_adj_658 : std_logic;
signal n5122 : std_logic;
signal \bluejay_data_inst.n14_cascade_\ : std_logic;
signal n5546 : std_logic;
signal \bluejay_data_inst.valid_o_N_155_cascade_\ : std_logic;
signal \bluejay_data_inst.n10\ : std_logic;
signal \bluejay_data_inst.n31_cascade_\ : std_logic;
signal \bluejay_data_inst.n4253_cascade_\ : std_logic;
signal \bluejay_data_inst.n1038_cascade_\ : std_logic;
signal \bluejay_data_inst.n31\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_7_N_122_5_cascade_\ : std_logic;
signal \DEBUG_3_c\ : std_logic;
signal \bluejay_data_inst.n11\ : std_logic;
signal \bluejay_data_inst.n9\ : std_logic;
signal \bluejay_data_inst.n4252\ : std_logic;
signal \bluejay_data_inst.n4_adj_648\ : std_logic;
signal \bluejay_data_inst.n3627_cascade_\ : std_logic;
signal \VALID_c\ : std_logic;
signal n5 : std_logic;
signal \bluejay_data_inst.n3631_cascade_\ : std_logic;
signal reset_all_w : std_logic;
signal \bluejay_data_inst.state_timeout_counter_7_N_122_5\ : std_logic;
signal \bluejay_data_inst.n4266\ : std_logic;
signal \bluejay_data_inst.n4_adj_652\ : std_logic;
signal \FIFO_D0_c_0\ : std_logic;
signal \DATA0_c_0\ : std_logic;
signal \DEBUG_6_c_22_c\ : std_logic;
signal \DEBUG_5_c\ : std_logic;
signal \r_SM_Main_2_adj_659\ : std_logic;
signal \pc_tx.n1\ : std_logic;
signal \bluejay_data_inst.h_counter_0\ : std_logic;
signal \bfn_17_7_0_\ : std_logic;
signal \bluejay_data_inst.h_counter_1\ : std_logic;
signal \bluejay_data_inst.n4858\ : std_logic;
signal \bluejay_data_inst.h_counter_2\ : std_logic;
signal \bluejay_data_inst.n4859\ : std_logic;
signal \bluejay_data_inst.h_counter_3\ : std_logic;
signal \bluejay_data_inst.n5547\ : std_logic;
signal \bluejay_data_inst.n4860\ : std_logic;
signal \bluejay_data_inst.h_counter_4\ : std_logic;
signal \bluejay_data_inst.n4861\ : std_logic;
signal \bluejay_data_inst.valid_o_N_155\ : std_logic;
signal \bluejay_data_inst.h_counter_5\ : std_logic;
signal \bluejay_data_inst.n5548\ : std_logic;
signal \bluejay_data_inst.n4862\ : std_logic;
signal \bluejay_data_inst.h_counter_6\ : std_logic;
signal \bluejay_data_inst.n4863\ : std_logic;
signal \bluejay_data_inst.n4864\ : std_logic;
signal \bluejay_data_inst.h_counter_7\ : std_logic;
signal n2555 : std_logic;
signal \bluejay_data_inst.n2693\ : std_logic;
signal \bfn_17_8_0_\ : std_logic;
signal \bluejay_data_inst.n5527\ : std_logic;
signal \bluejay_data_inst.n4816\ : std_logic;
signal \bluejay_data_inst.n51\ : std_logic;
signal \bluejay_data_inst.n4817\ : std_logic;
signal \bluejay_data_inst.n50\ : std_logic;
signal \bluejay_data_inst.n4818\ : std_logic;
signal \bluejay_data_inst.n4819\ : std_logic;
signal \bluejay_data_inst.n48\ : std_logic;
signal \bluejay_data_inst.n4820\ : std_logic;
signal \bluejay_data_inst.n4821\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \bluejay_data_inst.n4822\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_7_N_122_4_cascade_\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_7_N_122_4\ : std_logic;
signal \bluejay_data_inst.n8_cascade_\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_1\ : std_logic;
signal \bluejay_data_inst.n10_adj_654_cascade_\ : std_logic;
signal \bluejay_data_inst.n49\ : std_logic;
signal \bluejay_data_inst.n1394_cascade_\ : std_logic;
signal \bluejay_data_inst.n1039\ : std_logic;
signal \bluejay_data_inst.n4\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_4\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_3\ : std_logic;
signal \bluejay_data_inst.n14_adj_655\ : std_logic;
signal \bluejay_data_inst.n5544\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_7_N_122_7_cascade_\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_7_N_122_7\ : std_logic;
signal \bluejay_data_inst.n8_adj_640_cascade_\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_7\ : std_logic;
signal \bluejay_data_inst.n4_adj_641\ : std_logic;
signal \bluejay_data_inst.n5_adj_653\ : std_logic;
signal \bluejay_data_inst.n3602\ : std_logic;
signal n15 : std_logic;
signal \bluejay_data_inst.n1394\ : std_logic;
signal \bluejay_data_inst.n1133\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_5\ : std_logic;
signal \bluejay_data_inst.n4_adj_637\ : std_logic;
signal \FIFO_D4_c_4\ : std_logic;
signal \DATA4_c_4\ : std_logic;
signal \bluejay_data_inst.n5545\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_6\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_7_N_122_6_cascade_\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_7_N_122_6\ : std_logic;
signal \bluejay_data_inst.n8_adj_638_cascade_\ : std_logic;
signal \bluejay_data_inst.n4_adj_639\ : std_logic;
signal \bluejay_data_inst.n1054\ : std_logic;
signal \bluejay_data_inst.n5521\ : std_logic;
signal \bluejay_data_inst.n34\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_7_N_122_0_cascade_\ : std_logic;
signal \bluejay_data_inst.n8_adj_645_cascade_\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_7_N_122_0\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_7_N_122_2\ : std_logic;
signal n3_adj_669 : std_logic;
signal \bluejay_data_inst.n4260\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_2\ : std_logic;
signal \bluejay_data_inst.n4_adj_650\ : std_logic;
signal \bluejay_data_inst.state_timeout_counter_0\ : std_logic;
signal \bluejay_data_inst.n4_adj_636\ : std_logic;
signal \FIFO_D7_c_7\ : std_logic;
signal \DATA7_c_7\ : std_logic;
signal \FIFO_D17_c_17\ : std_logic;
signal \DATA17_c_17\ : std_logic;
signal \bluejay_data_inst.data_output_active_cmd\ : std_logic;
signal \FIFO_D2_c_2\ : std_logic;
signal \DATA2_c_2\ : std_logic;
signal get_next_word_cmd : std_logic;
signal \DEBUG_8_c\ : std_logic;
signal state_2 : std_logic;
signal \bluejay_data_inst.state_1\ : std_logic;
signal state_0 : std_logic;
signal \UPDATE_c\ : std_logic;
signal \bluejay_data_inst.n2096\ : std_logic;
signal \r_Rx_Data\ : std_logic;
signal n25_adj_662 : std_logic;
signal \bfn_23_5_0_\ : std_logic;
signal n24 : std_logic;
signal n4823 : std_logic;
signal n23 : std_logic;
signal n4824 : std_logic;
signal n22 : std_logic;
signal n4825 : std_logic;
signal n21 : std_logic;
signal n4826 : std_logic;
signal n20 : std_logic;
signal n4827 : std_logic;
signal n19 : std_logic;
signal n4828 : std_logic;
signal n18 : std_logic;
signal n4829 : std_logic;
signal n4830 : std_logic;
signal n17 : std_logic;
signal \bfn_23_6_0_\ : std_logic;
signal n16 : std_logic;
signal n4831 : std_logic;
signal n15_adj_663 : std_logic;
signal n4832 : std_logic;
signal n14 : std_logic;
signal n4833 : std_logic;
signal n13 : std_logic;
signal n4834 : std_logic;
signal n12 : std_logic;
signal n4835 : std_logic;
signal n11_adj_661 : std_logic;
signal n4836 : std_logic;
signal n10 : std_logic;
signal n4837 : std_logic;
signal n4838 : std_logic;
signal n9 : std_logic;
signal \bfn_23_7_0_\ : std_logic;
signal n8 : std_logic;
signal n4839 : std_logic;
signal n7 : std_logic;
signal n4840 : std_logic;
signal n6 : std_logic;
signal n4841 : std_logic;
signal n5_adj_665 : std_logic;
signal n4842 : std_logic;
signal n4_adj_664 : std_logic;
signal n4843 : std_logic;
signal n3 : std_logic;
signal n4844 : std_logic;
signal n2 : std_logic;
signal n4845 : std_logic;
signal n4846 : std_logic;
signal \bfn_23_8_0_\ : std_logic;
signal \DEBUG_0_c_24\ : std_logic;
signal \FR_RXF_c\ : std_logic;
signal \DEBUG_1_c\ : std_logic;
signal \GB_BUFFER_SLM_CLK_c_THRU_CO\ : std_logic;
signal \UART_RX_c\ : std_logic;
signal \pc_rx.r_Rx_Data_R\ : std_logic;
signal \SLM_CLK_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \FIFO_CLK_wire\ : std_logic;
signal \VALID_wire\ : std_logic;
signal \FIFO_D14_wire\ : std_logic;
signal \DATA30_wire\ : std_logic;
signal \DEBUG_9_wire\ : std_logic;
signal \FIFO_D8_wire\ : std_logic;
signal \DATA7_wire\ : std_logic;
signal \DEBUG_1_wire\ : std_logic;
signal \DATA4_wire\ : std_logic;
signal \FIFO_D26_wire\ : std_logic;
signal \DATA24_wire\ : std_logic;
signal \DTR_wire\ : std_logic;
signal \DATA29_wire\ : std_logic;
signal \FIFO_D16_wire\ : std_logic;
signal \FT_SIWU_wire\ : std_logic;
signal \DEBUG_6_wire\ : std_logic;
signal \DATA17_wire\ : std_logic;
signal \DATA21_wire\ : std_logic;
signal \DEBUG_5_wire\ : std_logic;
signal \DATA22_wire\ : std_logic;
signal \DSR_wire\ : std_logic;
signal \FT_WR_wire\ : std_logic;
signal \DATA26_wire\ : std_logic;
signal \FT_RD_wire\ : std_logic;
signal \DATA31_wire\ : std_logic;
signal \FIFO_D10_wire\ : std_logic;
signal \DATA5_wire\ : std_logic;
signal \INVERT_wire\ : std_logic;
signal \FIFO_D13_wire\ : std_logic;
signal \DEBUG_3_wire\ : std_logic;
signal \DATA8_wire\ : std_logic;
signal \DATA15_wire\ : std_logic;
signal \DATA20_wire\ : std_logic;
signal \DATA16_wire\ : std_logic;
signal \DATA28_wire\ : std_logic;
signal \FIFO_D23_wire\ : std_logic;
signal \CTS_wire\ : std_logic;
signal \SLM_CLK_wire\ : std_logic;
signal \FIFO_D20_wire\ : std_logic;
signal \FIFO_D19_wire\ : std_logic;
signal \FIFO_D7_wire\ : std_logic;
signal \UART_RX_wire\ : std_logic;
signal \FIFO_D6_wire\ : std_logic;
signal \DATA19_wire\ : std_logic;
signal \FIFO_D28_wire\ : std_logic;
signal \DATA14_wire\ : std_logic;
signal \DATA10_wire\ : std_logic;
signal \DATA6_wire\ : std_logic;
signal \FIFO_D11_wire\ : std_logic;
signal \FIFO_D3_wire\ : std_logic;
signal \RST_wire\ : std_logic;
signal \FIFO_D25_wire\ : std_logic;
signal \ICE_CDONE_wire\ : std_logic;
signal \SEN_wire\ : std_logic;
signal \DCD_wire\ : std_logic;
signal \FIFO_D9_wire\ : std_logic;
signal \DATA9_wire\ : std_logic;
signal \FIFO_D12_wire\ : std_logic;
signal \DATA27_wire\ : std_logic;
signal \DEBUG_0_wire\ : std_logic;
signal \DATA2_wire\ : std_logic;
signal \FIFO_D24_wire\ : std_logic;
signal \FIFO_D2_wire\ : std_logic;
signal \UART_TX_wire\ : std_logic;
signal \FIFO_D29_wire\ : std_logic;
signal \FIFO_D22_wire\ : std_logic;
signal \FIFO_D21_wire\ : std_logic;
signal \FR_RXF_wire\ : std_logic;
signal \DEBUG_8_wire\ : std_logic;
signal \FIFO_D15_wire\ : std_logic;
signal \DEBUG_2_wire\ : std_logic;
signal \DATA13_wire\ : std_logic;
signal \FIFO_D5_wire\ : std_logic;
signal \FIFO_D4_wire\ : std_logic;
signal \FIFO_D18_wire\ : std_logic;
signal \DATA23_wire\ : std_logic;
signal \FIFO_D30_wire\ : std_logic;
signal \DATA0_wire\ : std_logic;
signal \SYNC_wire\ : std_logic;
signal \SCK_wire\ : std_logic;
signal \UPDATE_wire\ : std_logic;
signal \DATA3_wire\ : std_logic;
signal \DATA18_wire\ : std_logic;
signal \DATA25_wire\ : std_logic;
signal \RESET_wire\ : std_logic;
signal \FIFO_D0_wire\ : std_logic;
signal \DATA12_wire\ : std_logic;
signal \FIFO_D31_wire\ : std_logic;
signal \SOUT_wire\ : std_logic;
signal \DATA11_wire\ : std_logic;
signal \DATA1_wire\ : std_logic;
signal \ICE_CREST_wire\ : std_logic;
signal \FIFO_D17_wire\ : std_logic;
signal \FIFO_D27_wire\ : std_logic;
signal \FIFO_D1_wire\ : std_logic;
signal \ICE_CLK_wire\ : std_logic;
signal \FT_OE_wire\ : std_logic;
signal \SDAT_wire\ : std_logic;

begin
    \FIFO_CLK_wire\ <= FIFO_CLK;
    VALID <= \VALID_wire\;
    \FIFO_D14_wire\ <= FIFO_D14;
    DATA30 <= \DATA30_wire\;
    DEBUG_9 <= \DEBUG_9_wire\;
    \FIFO_D8_wire\ <= FIFO_D8;
    DATA7 <= \DATA7_wire\;
    DEBUG_1 <= \DEBUG_1_wire\;
    DATA4 <= \DATA4_wire\;
    \FIFO_D26_wire\ <= FIFO_D26;
    DATA24 <= \DATA24_wire\;
    DTR <= \DTR_wire\;
    DATA29 <= \DATA29_wire\;
    \FIFO_D16_wire\ <= FIFO_D16;
    FT_SIWU <= \FT_SIWU_wire\;
    DEBUG_6 <= \DEBUG_6_wire\;
    DATA17 <= \DATA17_wire\;
    DATA21 <= \DATA21_wire\;
    DEBUG_5 <= \DEBUG_5_wire\;
    DATA22 <= \DATA22_wire\;
    DSR <= \DSR_wire\;
    FT_WR <= \FT_WR_wire\;
    DATA26 <= \DATA26_wire\;
    FT_RD <= \FT_RD_wire\;
    DATA31 <= \DATA31_wire\;
    \FIFO_D10_wire\ <= FIFO_D10;
    DATA5 <= \DATA5_wire\;
    INVERT <= \INVERT_wire\;
    \FIFO_D13_wire\ <= FIFO_D13;
    DEBUG_3 <= \DEBUG_3_wire\;
    DATA8 <= \DATA8_wire\;
    DATA15 <= \DATA15_wire\;
    DATA20 <= \DATA20_wire\;
    DATA16 <= \DATA16_wire\;
    DATA28 <= \DATA28_wire\;
    \FIFO_D23_wire\ <= FIFO_D23;
    CTS <= \CTS_wire\;
    SLM_CLK <= \SLM_CLK_wire\;
    \FIFO_D20_wire\ <= FIFO_D20;
    \FIFO_D19_wire\ <= FIFO_D19;
    \FIFO_D7_wire\ <= FIFO_D7;
    \UART_RX_wire\ <= UART_RX;
    \FIFO_D6_wire\ <= FIFO_D6;
    DATA19 <= \DATA19_wire\;
    \FIFO_D28_wire\ <= FIFO_D28;
    DATA14 <= \DATA14_wire\;
    DATA10 <= \DATA10_wire\;
    DATA6 <= \DATA6_wire\;
    \FIFO_D11_wire\ <= FIFO_D11;
    \FIFO_D3_wire\ <= FIFO_D3;
    RST <= \RST_wire\;
    \FIFO_D25_wire\ <= FIFO_D25;
    ICE_CDONE <= \ICE_CDONE_wire\;
    SEN <= \SEN_wire\;
    DCD <= \DCD_wire\;
    \FIFO_D9_wire\ <= FIFO_D9;
    DATA9 <= \DATA9_wire\;
    \FIFO_D12_wire\ <= FIFO_D12;
    DATA27 <= \DATA27_wire\;
    DEBUG_0 <= \DEBUG_0_wire\;
    DATA2 <= \DATA2_wire\;
    \FIFO_D24_wire\ <= FIFO_D24;
    \FIFO_D2_wire\ <= FIFO_D2;
    UART_TX <= \UART_TX_wire\;
    \FIFO_D29_wire\ <= FIFO_D29;
    \FIFO_D22_wire\ <= FIFO_D22;
    \FIFO_D21_wire\ <= FIFO_D21;
    \FR_RXF_wire\ <= FR_RXF;
    DEBUG_8 <= \DEBUG_8_wire\;
    \FIFO_D15_wire\ <= FIFO_D15;
    DEBUG_2 <= \DEBUG_2_wire\;
    DATA13 <= \DATA13_wire\;
    \FIFO_D5_wire\ <= FIFO_D5;
    \FIFO_D4_wire\ <= FIFO_D4;
    \FIFO_D18_wire\ <= FIFO_D18;
    DATA23 <= \DATA23_wire\;
    \FIFO_D30_wire\ <= FIFO_D30;
    DATA0 <= \DATA0_wire\;
    SYNC <= \SYNC_wire\;
    SCK <= \SCK_wire\;
    UPDATE <= \UPDATE_wire\;
    DATA3 <= \DATA3_wire\;
    DATA18 <= \DATA18_wire\;
    DATA25 <= \DATA25_wire\;
    RESET <= \RESET_wire\;
    \FIFO_D0_wire\ <= FIFO_D0;
    DATA12 <= \DATA12_wire\;
    \FIFO_D31_wire\ <= FIFO_D31;
    \SOUT_wire\ <= SOUT;
    DATA11 <= \DATA11_wire\;
    DATA1 <= \DATA1_wire\;
    ICE_CREST <= \ICE_CREST_wire\;
    \FIFO_D17_wire\ <= FIFO_D17;
    \FIFO_D27_wire\ <= FIFO_D27;
    \FIFO_D1_wire\ <= FIFO_D1;
    ICE_CLK <= \ICE_CLK_wire\;
    FT_OE <= \FT_OE_wire\;
    SDAT <= \SDAT_wire\;

    \FIFO_CLK_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__20522\,
            GLOBALBUFFEROUTPUT => \SLM_CLK_c\
        );

    \FIFO_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20524\,
            DIN => \N__20523\,
            DOUT => \N__20522\,
            PACKAGEPIN => \FIFO_CLK_wire\
        );

    \FIFO_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20524\,
            PADOUT => \N__20523\,
            PADIN => \N__20522\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VALID_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20513\,
            DIN => \N__20512\,
            DOUT => \N__20511\,
            PACKAGEPIN => \VALID_wire\
        );

    \VALID_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20513\,
            PADOUT => \N__20512\,
            PADIN => \N__20511\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__15931\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D14_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20504\,
            DIN => \N__20503\,
            DOUT => \N__20502\,
            PACKAGEPIN => \FIFO_D14_wire\
        );

    \FIFO_D14_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20504\,
            PADOUT => \N__20503\,
            PADIN => \N__20502\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D14_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA30_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20495\,
            DIN => \N__20494\,
            DOUT => \N__20493\,
            PACKAGEPIN => \DATA30_wire\
        );

    \DATA30_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20495\,
            PADOUT => \N__20494\,
            PADIN => \N__20493\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7465\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_9_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20486\,
            DIN => \N__20485\,
            DOUT => \N__20484\,
            PACKAGEPIN => \DEBUG_9_wire\
        );

    \DEBUG_9_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20486\,
            PADOUT => \N__20485\,
            PADIN => \N__20484\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10839\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D8_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20477\,
            DIN => \N__20476\,
            DOUT => \N__20475\,
            PACKAGEPIN => \FIFO_D8_wire\
        );

    \FIFO_D8_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20477\,
            PADOUT => \N__20476\,
            PADIN => \N__20475\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D8_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA7_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20468\,
            DIN => \N__20467\,
            DOUT => \N__20466\,
            PACKAGEPIN => \DATA7_wire\
        );

    \DATA7_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20468\,
            PADOUT => \N__20467\,
            PADIN => \N__20466\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17608\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20459\,
            DIN => \N__20458\,
            DOUT => \N__20457\,
            PACKAGEPIN => \DEBUG_1_wire\
        );

    \DEBUG_1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20459\,
            PADOUT => \N__20458\,
            PADIN => \N__20457\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19459\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA4_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20450\,
            DIN => \N__20449\,
            DOUT => \N__20448\,
            PACKAGEPIN => \DATA4_wire\
        );

    \DATA4_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20450\,
            PADOUT => \N__20449\,
            PADIN => \N__20448\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17344\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D26_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20441\,
            DIN => \N__20440\,
            DOUT => \N__20439\,
            PACKAGEPIN => \FIFO_D26_wire\
        );

    \FIFO_D26_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20441\,
            PADOUT => \N__20440\,
            PADIN => \N__20439\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D26_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA24_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20432\,
            DIN => \N__20431\,
            DOUT => \N__20430\,
            PACKAGEPIN => \DATA24_wire\
        );

    \DATA24_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20432\,
            PADOUT => \N__20431\,
            PADIN => \N__20430\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12580\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DTR_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20423\,
            DIN => \N__20422\,
            DOUT => \N__20421\,
            PACKAGEPIN => \DTR_wire\
        );

    \DTR_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20423\,
            PADOUT => \N__20422\,
            PADIN => \N__20421\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA29_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20414\,
            DIN => \N__20413\,
            DOUT => \N__20412\,
            PACKAGEPIN => \DATA29_wire\
        );

    \DATA29_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20414\,
            PADOUT => \N__20413\,
            PADIN => \N__20412\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8137\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D16_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20405\,
            DIN => \N__20404\,
            DOUT => \N__20403\,
            PACKAGEPIN => \FIFO_D16_wire\
        );

    \FIFO_D16_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20405\,
            PADOUT => \N__20404\,
            PADIN => \N__20403\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D16_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FT_SIWU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20396\,
            DIN => \N__20395\,
            DOUT => \N__20394\,
            PACKAGEPIN => \FT_SIWU_wire\
        );

    \FT_SIWU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20396\,
            PADOUT => \N__20395\,
            PADIN => \N__20394\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17115\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_6_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20387\,
            DIN => \N__20386\,
            DOUT => \N__20385\,
            PACKAGEPIN => \DEBUG_6_wire\
        );

    \DEBUG_6_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20387\,
            PADOUT => \N__20386\,
            PADIN => \N__20385\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16249\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA17_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20378\,
            DIN => \N__20377\,
            DOUT => \N__20376\,
            PACKAGEPIN => \DATA17_wire\
        );

    \DATA17_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20378\,
            PADOUT => \N__20377\,
            PADIN => \N__20376\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18991\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA21_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20369\,
            DIN => \N__20368\,
            DOUT => \N__20367\,
            PACKAGEPIN => \DATA21_wire\
        );

    \DATA21_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20369\,
            PADOUT => \N__20368\,
            PADIN => \N__20367\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13189\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_5_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20360\,
            DIN => \N__20359\,
            DOUT => \N__20358\,
            PACKAGEPIN => \DEBUG_5_wire\
        );

    \DEBUG_5_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20360\,
            PADOUT => \N__20359\,
            PADIN => \N__20358\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16200\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA22_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20351\,
            DIN => \N__20350\,
            DOUT => \N__20349\,
            PACKAGEPIN => \DATA22_wire\
        );

    \DATA22_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20351\,
            PADOUT => \N__20350\,
            PADIN => \N__20349\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16210\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DSR_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20342\,
            DIN => \N__20341\,
            DOUT => \N__20340\,
            PACKAGEPIN => \DSR_wire\
        );

    \DSR_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20342\,
            PADOUT => \N__20341\,
            PADIN => \N__20340\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FT_WR_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20333\,
            DIN => \N__20332\,
            DOUT => \N__20331\,
            PACKAGEPIN => \FT_WR_wire\
        );

    \FT_WR_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20333\,
            PADOUT => \N__20332\,
            PADIN => \N__20331\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17119\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA26_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20324\,
            DIN => \N__20323\,
            DOUT => \N__20322\,
            PACKAGEPIN => \DATA26_wire\
        );

    \DATA26_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20324\,
            PADOUT => \N__20323\,
            PADIN => \N__20322\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10339\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FT_RD_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20315\,
            DIN => \N__20314\,
            DOUT => \N__20313\,
            PACKAGEPIN => \FT_RD_wire\
        );

    \FT_RD_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20315\,
            PADOUT => \N__20314\,
            PADIN => \N__20313\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7584\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA31_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20306\,
            DIN => \N__20305\,
            DOUT => \N__20304\,
            PACKAGEPIN => \DATA31_wire\
        );

    \DATA31_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20306\,
            PADOUT => \N__20305\,
            PADIN => \N__20304\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7687\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D10_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20297\,
            DIN => \N__20296\,
            DOUT => \N__20295\,
            PACKAGEPIN => \FIFO_D10_wire\
        );

    \FIFO_D10_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20297\,
            PADOUT => \N__20296\,
            PADIN => \N__20295\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D10_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA5_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20288\,
            DIN => \N__20287\,
            DOUT => \N__20286\,
            PACKAGEPIN => \DATA5_wire\
        );

    \DATA5_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20288\,
            PADOUT => \N__20287\,
            PADIN => \N__20286\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12547\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \INVERT_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20279\,
            DIN => \N__20278\,
            DOUT => \N__20277\,
            PACKAGEPIN => \INVERT_wire\
        );

    \INVERT_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20279\,
            PADOUT => \N__20278\,
            PADIN => \N__20277\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D13_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20270\,
            DIN => \N__20269\,
            DOUT => \N__20268\,
            PACKAGEPIN => \FIFO_D13_wire\
        );

    \FIFO_D13_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20270\,
            PADOUT => \N__20269\,
            PADIN => \N__20268\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D13_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20261\,
            DIN => \N__20260\,
            DOUT => \N__20259\,
            PACKAGEPIN => \DEBUG_3_wire\
        );

    \DEBUG_3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20261\,
            PADOUT => \N__20260\,
            PADIN => \N__20259\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16003\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA8_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20252\,
            DIN => \N__20251\,
            DOUT => \N__20250\,
            PACKAGEPIN => \DATA8_wire\
        );

    \DATA8_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20252\,
            PADOUT => \N__20251\,
            PADIN => \N__20250\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9631\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA15_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20243\,
            DIN => \N__20242\,
            DOUT => \N__20241\,
            PACKAGEPIN => \DATA15_wire\
        );

    \DATA15_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20243\,
            PADOUT => \N__20242\,
            PADIN => \N__20241\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10786\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA20_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20234\,
            DIN => \N__20233\,
            DOUT => \N__20232\,
            PACKAGEPIN => \DATA20_wire\
        );

    \DATA20_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20234\,
            PADOUT => \N__20233\,
            PADIN => \N__20232\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11512\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA16_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20225\,
            DIN => \N__20224\,
            DOUT => \N__20223\,
            PACKAGEPIN => \DATA16_wire\
        );

    \DATA16_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20225\,
            PADOUT => \N__20224\,
            PADIN => \N__20223\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14044\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA28_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20216\,
            DIN => \N__20215\,
            DOUT => \N__20214\,
            PACKAGEPIN => \DATA28_wire\
        );

    \DATA28_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20216\,
            PADOUT => \N__20215\,
            PADIN => \N__20214\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7834\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D23_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20207\,
            DIN => \N__20206\,
            DOUT => \N__20205\,
            PACKAGEPIN => \FIFO_D23_wire\
        );

    \FIFO_D23_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20207\,
            PADOUT => \N__20206\,
            PADIN => \N__20205\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D23_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CTS_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20198\,
            DIN => \N__20197\,
            DOUT => \N__20196\,
            PACKAGEPIN => \CTS_wire\
        );

    \CTS_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20198\,
            PADOUT => \N__20197\,
            PADIN => \N__20196\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SLM_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20189\,
            DIN => \N__20188\,
            DOUT => \N__20187\,
            PACKAGEPIN => \SLM_CLK_wire\
        );

    \SLM_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20189\,
            PADOUT => \N__20188\,
            PADIN => \N__20187\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19447\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D20_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20180\,
            DIN => \N__20179\,
            DOUT => \N__20178\,
            PACKAGEPIN => \FIFO_D20_wire\
        );

    \FIFO_D20_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20180\,
            PADOUT => \N__20179\,
            PADIN => \N__20178\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D20_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D19_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20171\,
            DIN => \N__20170\,
            DOUT => \N__20169\,
            PACKAGEPIN => \FIFO_D19_wire\
        );

    \FIFO_D19_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20171\,
            PADOUT => \N__20170\,
            PADIN => \N__20169\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D19_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D7_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20162\,
            DIN => \N__20161\,
            DOUT => \N__20160\,
            PACKAGEPIN => \FIFO_D7_wire\
        );

    \FIFO_D7_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20162\,
            PADOUT => \N__20161\,
            PADIN => \N__20160\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D7_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UART_RX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20153\,
            DIN => \N__20152\,
            DOUT => \N__20151\,
            PACKAGEPIN => \UART_RX_wire\
        );

    \UART_RX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20153\,
            PADOUT => \N__20152\,
            PADIN => \N__20151\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \UART_RX_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D6_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20144\,
            DIN => \N__20143\,
            DOUT => \N__20142\,
            PACKAGEPIN => \FIFO_D6_wire\
        );

    \FIFO_D6_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20144\,
            PADOUT => \N__20143\,
            PADIN => \N__20142\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D6_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA19_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20135\,
            DIN => \N__20134\,
            DOUT => \N__20133\,
            PACKAGEPIN => \DATA19_wire\
        );

    \DATA19_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20135\,
            PADOUT => \N__20134\,
            PADIN => \N__20133\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7549\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D28_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20126\,
            DIN => \N__20125\,
            DOUT => \N__20124\,
            PACKAGEPIN => \FIFO_D28_wire\
        );

    \FIFO_D28_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20126\,
            PADOUT => \N__20125\,
            PADIN => \N__20124\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D28_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA14_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20117\,
            DIN => \N__20116\,
            DOUT => \N__20115\,
            PACKAGEPIN => \DATA14_wire\
        );

    \DATA14_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20117\,
            PADOUT => \N__20116\,
            PADIN => \N__20115\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7504\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA10_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20108\,
            DIN => \N__20107\,
            DOUT => \N__20106\,
            PACKAGEPIN => \DATA10_wire\
        );

    \DATA10_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20108\,
            PADOUT => \N__20107\,
            PADIN => \N__20106\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14128\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA6_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20099\,
            DIN => \N__20098\,
            DOUT => \N__20097\,
            PACKAGEPIN => \DATA6_wire\
        );

    \DATA6_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20099\,
            PADOUT => \N__20098\,
            PADIN => \N__20097\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12514\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D11_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20090\,
            DIN => \N__20089\,
            DOUT => \N__20088\,
            PACKAGEPIN => \FIFO_D11_wire\
        );

    \FIFO_D11_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20090\,
            PADOUT => \N__20089\,
            PADIN => \N__20088\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D11_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20081\,
            DIN => \N__20080\,
            DOUT => \N__20079\,
            PACKAGEPIN => \FIFO_D3_wire\
        );

    \FIFO_D3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20081\,
            PADOUT => \N__20080\,
            PADIN => \N__20079\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D3_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RST_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20072\,
            DIN => \N__20071\,
            DOUT => \N__20070\,
            PACKAGEPIN => \RST_wire\
        );

    \RST_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20072\,
            PADOUT => \N__20071\,
            PADIN => \N__20070\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D25_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20063\,
            DIN => \N__20062\,
            DOUT => \N__20061\,
            PACKAGEPIN => \FIFO_D25_wire\
        );

    \FIFO_D25_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20063\,
            PADOUT => \N__20062\,
            PADIN => \N__20061\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D25_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ICE_CDONE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20054\,
            DIN => \N__20053\,
            DOUT => \N__20052\,
            PACKAGEPIN => \ICE_CDONE_wire\
        );

    \ICE_CDONE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20054\,
            PADOUT => \N__20053\,
            PADIN => \N__20052\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SEN_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20045\,
            DIN => \N__20044\,
            DOUT => \N__20043\,
            PACKAGEPIN => \SEN_wire\
        );

    \SEN_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20045\,
            PADOUT => \N__20044\,
            PADIN => \N__20043\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8221\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DCD_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20036\,
            DIN => \N__20035\,
            DOUT => \N__20034\,
            PACKAGEPIN => \DCD_wire\
        );

    \DCD_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20036\,
            PADOUT => \N__20035\,
            PADIN => \N__20034\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D9_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20027\,
            DIN => \N__20026\,
            DOUT => \N__20025\,
            PACKAGEPIN => \FIFO_D9_wire\
        );

    \FIFO_D9_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20027\,
            PADOUT => \N__20026\,
            PADIN => \N__20025\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D9_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA9_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20018\,
            DIN => \N__20017\,
            DOUT => \N__20016\,
            PACKAGEPIN => \DATA9_wire\
        );

    \DATA9_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20018\,
            PADOUT => \N__20017\,
            PADIN => \N__20016\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14089\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D12_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20009\,
            DIN => \N__20008\,
            DOUT => \N__20007\,
            PACKAGEPIN => \FIFO_D12_wire\
        );

    \FIFO_D12_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20009\,
            PADOUT => \N__20008\,
            PADIN => \N__20007\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D12_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA27_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20000\,
            DIN => \N__19999\,
            DOUT => \N__19998\,
            PACKAGEPIN => \DATA27_wire\
        );

    \DATA27_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20000\,
            PADOUT => \N__19999\,
            PADIN => \N__19998\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11551\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_0_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19991\,
            DIN => \N__19990\,
            DOUT => \N__19989\,
            PACKAGEPIN => \DEBUG_0_wire\
        );

    \DEBUG_0_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19991\,
            PADOUT => \N__19990\,
            PADIN => \N__19989\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19591\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19982\,
            DIN => \N__19981\,
            DOUT => \N__19980\,
            PACKAGEPIN => \DATA2_wire\
        );

    \DATA2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19982\,
            PADOUT => \N__19981\,
            PADIN => \N__19980\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18679\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D24_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19973\,
            DIN => \N__19972\,
            DOUT => \N__19971\,
            PACKAGEPIN => \FIFO_D24_wire\
        );

    \FIFO_D24_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19973\,
            PADOUT => \N__19972\,
            PADIN => \N__19971\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D24_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19964\,
            DIN => \N__19963\,
            DOUT => \N__19962\,
            PACKAGEPIN => \FIFO_D2_wire\
        );

    \FIFO_D2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19964\,
            PADOUT => \N__19963\,
            PADIN => \N__19962\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D2_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UART_TX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19955\,
            DIN => \N__19954\,
            DOUT => \N__19953\,
            PACKAGEPIN => \UART_TX_wire\
        );

    \UART_TX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19955\,
            PADOUT => \N__19954\,
            PADIN => \N__19953\,
            CLOCKENABLE => \N__16096\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9100\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__19404\
        );

    \FIFO_D29_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19946\,
            DIN => \N__19945\,
            DOUT => \N__19944\,
            PACKAGEPIN => \FIFO_D29_wire\
        );

    \FIFO_D29_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19946\,
            PADOUT => \N__19945\,
            PADIN => \N__19944\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D29_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_6_c_22_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19937\,
            DIN => \N__19936\,
            DOUT => \N__19935\,
            PACKAGEPIN => \FIFO_D22_wire\
        );

    \DEBUG_6_c_22_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19937\,
            PADOUT => \N__19936\,
            PADIN => \N__19935\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_6_c_22_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D21_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19928\,
            DIN => \N__19927\,
            DOUT => \N__19926\,
            PACKAGEPIN => \FIFO_D21_wire\
        );

    \FIFO_D21_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19928\,
            PADOUT => \N__19927\,
            PADIN => \N__19926\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D21_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FR_RXF_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19919\,
            DIN => \N__19918\,
            DOUT => \N__19917\,
            PACKAGEPIN => \FR_RXF_wire\
        );

    \FR_RXF_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19919\,
            PADOUT => \N__19918\,
            PADIN => \N__19917\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FR_RXF_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_8_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19910\,
            DIN => \N__19909\,
            DOUT => \N__19908\,
            PACKAGEPIN => \DEBUG_8_wire\
        );

    \DEBUG_8_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19910\,
            PADOUT => \N__19909\,
            PADIN => \N__19908\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18622\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D15_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19901\,
            DIN => \N__19900\,
            DOUT => \N__19899\,
            PACKAGEPIN => \FIFO_D15_wire\
        );

    \FIFO_D15_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19901\,
            PADOUT => \N__19900\,
            PADIN => \N__19899\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D15_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19892\,
            DIN => \N__19891\,
            DOUT => \N__19890\,
            PACKAGEPIN => \DEBUG_2_wire\
        );

    \DEBUG_2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19892\,
            PADOUT => \N__19891\,
            PADIN => \N__19890\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA13_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19883\,
            DIN => \N__19882\,
            DOUT => \N__19881\,
            PACKAGEPIN => \DATA13_wire\
        );

    \DATA13_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19883\,
            PADOUT => \N__19882\,
            PADIN => \N__19881\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11467\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D5_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19874\,
            DIN => \N__19873\,
            DOUT => \N__19872\,
            PACKAGEPIN => \FIFO_D5_wire\
        );

    \FIFO_D5_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19874\,
            PADOUT => \N__19873\,
            PADIN => \N__19872\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D5_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D4_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19865\,
            DIN => \N__19864\,
            DOUT => \N__19863\,
            PACKAGEPIN => \FIFO_D4_wire\
        );

    \FIFO_D4_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19865\,
            PADOUT => \N__19864\,
            PADIN => \N__19863\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D4_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D18_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19856\,
            DIN => \N__19855\,
            DOUT => \N__19854\,
            PACKAGEPIN => \FIFO_D18_wire\
        );

    \FIFO_D18_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19856\,
            PADOUT => \N__19855\,
            PADIN => \N__19854\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D18_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA23_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19847\,
            DIN => \N__19846\,
            DOUT => \N__19845\,
            PACKAGEPIN => \DATA23_wire\
        );

    \DATA23_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19847\,
            PADOUT => \N__19846\,
            PADIN => \N__19845\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7783\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D30_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19838\,
            DIN => \N__19837\,
            DOUT => \N__19836\,
            PACKAGEPIN => \FIFO_D30_wire\
        );

    \FIFO_D30_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19838\,
            PADOUT => \N__19837\,
            PADIN => \N__19836\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D30_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA0_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19829\,
            DIN => \N__19828\,
            DOUT => \N__19827\,
            PACKAGEPIN => \DATA0_wire\
        );

    \DATA0_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19829\,
            PADOUT => \N__19828\,
            PADIN => \N__19827\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16270\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19820\,
            DIN => \N__19819\,
            DOUT => \N__19818\,
            PACKAGEPIN => \SYNC_wire\
        );

    \SYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19820\,
            PADOUT => \N__19819\,
            PADIN => \N__19818\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SCK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19811\,
            DIN => \N__19810\,
            DOUT => \N__19809\,
            PACKAGEPIN => \SCK_wire\
        );

    \SCK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19811\,
            PADOUT => \N__19810\,
            PADIN => \N__19809\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7816\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UPDATE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19802\,
            DIN => \N__19801\,
            DOUT => \N__19800\,
            PACKAGEPIN => \UPDATE_wire\
        );

    \UPDATE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19802\,
            PADOUT => \N__19801\,
            PADIN => \N__19800\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18103\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19793\,
            DIN => \N__19792\,
            DOUT => \N__19791\,
            PACKAGEPIN => \DATA3_wire\
        );

    \DATA3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19793\,
            PADOUT => \N__19792\,
            PADIN => \N__19791\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__15148\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA18_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19784\,
            DIN => \N__19783\,
            DOUT => \N__19782\,
            PACKAGEPIN => \DATA18_wire\
        );

    \DATA18_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19784\,
            PADOUT => \N__19783\,
            PADIN => \N__19782\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8785\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA25_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19775\,
            DIN => \N__19774\,
            DOUT => \N__19773\,
            PACKAGEPIN => \DATA25_wire\
        );

    \DATA25_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19775\,
            PADOUT => \N__19774\,
            PADIN => \N__19773\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8173\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESET_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19766\,
            DIN => \N__19765\,
            DOUT => \N__19764\,
            PACKAGEPIN => \RESET_wire\
        );

    \RESET_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19766\,
            PADOUT => \N__19765\,
            PADIN => \N__19764\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11401\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D0_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19757\,
            DIN => \N__19756\,
            DOUT => \N__19755\,
            PACKAGEPIN => \FIFO_D0_wire\
        );

    \FIFO_D0_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19757\,
            PADOUT => \N__19756\,
            PADIN => \N__19755\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D0_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA12_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19748\,
            DIN => \N__19747\,
            DOUT => \N__19746\,
            PACKAGEPIN => \DATA12_wire\
        );

    \DATA12_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19748\,
            PADOUT => \N__19747\,
            PADIN => \N__19746\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__15109\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D31_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19739\,
            DIN => \N__19738\,
            DOUT => \N__19737\,
            PACKAGEPIN => \FIFO_D31_wire\
        );

    \FIFO_D31_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19739\,
            PADOUT => \N__19738\,
            PADIN => \N__19737\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D31_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SOUT_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19730\,
            DIN => \N__19729\,
            DOUT => \N__19728\,
            PACKAGEPIN => \SOUT_wire\
        );

    \SOUT_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19730\,
            PADOUT => \N__19729\,
            PADIN => \N__19728\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SOUT_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA11_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19721\,
            DIN => \N__19720\,
            DOUT => \N__19719\,
            PACKAGEPIN => \DATA11_wire\
        );

    \DATA11_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19721\,
            PADOUT => \N__19720\,
            PADIN => \N__19719\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7648\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19712\,
            DIN => \N__19711\,
            DOUT => \N__19710\,
            PACKAGEPIN => \DATA1_wire\
        );

    \DATA1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19712\,
            PADOUT => \N__19711\,
            PADIN => \N__19710\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13231\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ICE_CREST_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19703\,
            DIN => \N__19702\,
            DOUT => \N__19701\,
            PACKAGEPIN => \ICE_CREST_wire\
        );

    \ICE_CREST_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19703\,
            PADOUT => \N__19702\,
            PADIN => \N__19701\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D17_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19694\,
            DIN => \N__19693\,
            DOUT => \N__19692\,
            PACKAGEPIN => \FIFO_D17_wire\
        );

    \FIFO_D17_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19694\,
            PADOUT => \N__19693\,
            PADIN => \N__19692\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D17_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D27_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19685\,
            DIN => \N__19684\,
            DOUT => \N__19683\,
            PACKAGEPIN => \FIFO_D27_wire\
        );

    \FIFO_D27_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19685\,
            PADOUT => \N__19684\,
            PADIN => \N__19683\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D27_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19676\,
            DIN => \N__19675\,
            DOUT => \N__19674\,
            PACKAGEPIN => \FIFO_D1_wire\
        );

    \FIFO_D1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19676\,
            PADOUT => \N__19675\,
            PADIN => \N__19674\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \FIFO_D1_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ICE_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19667\,
            DIN => \N__19666\,
            DOUT => \N__19665\,
            PACKAGEPIN => \ICE_CLK_wire\
        );

    \ICE_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19667\,
            PADOUT => \N__19666\,
            PADIN => \N__19665\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FT_OE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19658\,
            DIN => \N__19657\,
            DOUT => \N__19656\,
            PACKAGEPIN => \FT_OE_wire\
        );

    \FT_OE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19658\,
            PADOUT => \N__19657\,
            PADIN => \N__19656\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7588\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SDAT_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19649\,
            DIN => \N__19648\,
            DOUT => \N__19647\,
            PACKAGEPIN => \SDAT_wire\
        );

    \SDAT_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19649\,
            PADOUT => \N__19648\,
            PADIN => \N__19647\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10843\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__4692\ : InMux
    port map (
            O => \N__19630\,
            I => \N__19627\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__19627\,
            I => n5_adj_665
        );

    \I__4690\ : InMux
    port map (
            O => \N__19624\,
            I => n4842
        );

    \I__4689\ : InMux
    port map (
            O => \N__19621\,
            I => \N__19618\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__19618\,
            I => n4_adj_664
        );

    \I__4687\ : InMux
    port map (
            O => \N__19615\,
            I => n4843
        );

    \I__4686\ : InMux
    port map (
            O => \N__19612\,
            I => \N__19609\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__19609\,
            I => n3
        );

    \I__4684\ : InMux
    port map (
            O => \N__19606\,
            I => n4844
        );

    \I__4683\ : InMux
    port map (
            O => \N__19603\,
            I => \N__19600\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__19600\,
            I => n2
        );

    \I__4681\ : InMux
    port map (
            O => \N__19597\,
            I => n4845
        );

    \I__4680\ : InMux
    port map (
            O => \N__19594\,
            I => \bfn_23_8_0_\
        );

    \I__4679\ : IoInMux
    port map (
            O => \N__19591\,
            I => \N__19588\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__19588\,
            I => \N__19585\
        );

    \I__4677\ : Span4Mux_s2_h
    port map (
            O => \N__19585\,
            I => \N__19582\
        );

    \I__4676\ : Span4Mux_v
    port map (
            O => \N__19582\,
            I => \N__19579\
        );

    \I__4675\ : Span4Mux_v
    port map (
            O => \N__19579\,
            I => \N__19575\
        );

    \I__4674\ : InMux
    port map (
            O => \N__19578\,
            I => \N__19572\
        );

    \I__4673\ : Odrv4
    port map (
            O => \N__19575\,
            I => \DEBUG_0_c_24\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__19572\,
            I => \DEBUG_0_c_24\
        );

    \I__4671\ : InMux
    port map (
            O => \N__19567\,
            I => \N__19562\
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__19566\,
            I => \N__19557\
        );

    \I__4669\ : InMux
    port map (
            O => \N__19565\,
            I => \N__19553\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__19562\,
            I => \N__19550\
        );

    \I__4667\ : InMux
    port map (
            O => \N__19561\,
            I => \N__19547\
        );

    \I__4666\ : InMux
    port map (
            O => \N__19560\,
            I => \N__19544\
        );

    \I__4665\ : InMux
    port map (
            O => \N__19557\,
            I => \N__19541\
        );

    \I__4664\ : CascadeMux
    port map (
            O => \N__19556\,
            I => \N__19538\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__19553\,
            I => \N__19535\
        );

    \I__4662\ : Span4Mux_v
    port map (
            O => \N__19550\,
            I => \N__19532\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__19547\,
            I => \N__19527\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__19544\,
            I => \N__19527\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__19541\,
            I => \N__19524\
        );

    \I__4658\ : InMux
    port map (
            O => \N__19538\,
            I => \N__19521\
        );

    \I__4657\ : Span4Mux_v
    port map (
            O => \N__19535\,
            I => \N__19518\
        );

    \I__4656\ : Span4Mux_h
    port map (
            O => \N__19532\,
            I => \N__19513\
        );

    \I__4655\ : Span4Mux_v
    port map (
            O => \N__19527\,
            I => \N__19513\
        );

    \I__4654\ : Span4Mux_v
    port map (
            O => \N__19524\,
            I => \N__19508\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__19521\,
            I => \N__19508\
        );

    \I__4652\ : Sp12to4
    port map (
            O => \N__19518\,
            I => \N__19504\
        );

    \I__4651\ : Span4Mux_h
    port map (
            O => \N__19513\,
            I => \N__19501\
        );

    \I__4650\ : Span4Mux_h
    port map (
            O => \N__19508\,
            I => \N__19498\
        );

    \I__4649\ : InMux
    port map (
            O => \N__19507\,
            I => \N__19495\
        );

    \I__4648\ : Span12Mux_h
    port map (
            O => \N__19504\,
            I => \N__19490\
        );

    \I__4647\ : Sp12to4
    port map (
            O => \N__19501\,
            I => \N__19490\
        );

    \I__4646\ : Span4Mux_h
    port map (
            O => \N__19498\,
            I => \N__19487\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__19495\,
            I => \N__19484\
        );

    \I__4644\ : Span12Mux_h
    port map (
            O => \N__19490\,
            I => \N__19481\
        );

    \I__4643\ : Sp12to4
    port map (
            O => \N__19487\,
            I => \N__19478\
        );

    \I__4642\ : Span4Mux_v
    port map (
            O => \N__19484\,
            I => \N__19475\
        );

    \I__4641\ : Span12Mux_v
    port map (
            O => \N__19481\,
            I => \N__19472\
        );

    \I__4640\ : Span12Mux_v
    port map (
            O => \N__19478\,
            I => \N__19469\
        );

    \I__4639\ : Span4Mux_h
    port map (
            O => \N__19475\,
            I => \N__19466\
        );

    \I__4638\ : Odrv12
    port map (
            O => \N__19472\,
            I => \FR_RXF_c\
        );

    \I__4637\ : Odrv12
    port map (
            O => \N__19469\,
            I => \FR_RXF_c\
        );

    \I__4636\ : Odrv4
    port map (
            O => \N__19466\,
            I => \FR_RXF_c\
        );

    \I__4635\ : IoInMux
    port map (
            O => \N__19459\,
            I => \N__19456\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__19456\,
            I => \N__19453\
        );

    \I__4633\ : Span12Mux_s5_h
    port map (
            O => \N__19453\,
            I => \N__19450\
        );

    \I__4632\ : Odrv12
    port map (
            O => \N__19450\,
            I => \DEBUG_1_c\
        );

    \I__4631\ : IoInMux
    port map (
            O => \N__19447\,
            I => \N__19444\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__19444\,
            I => \N__19441\
        );

    \I__4629\ : Span4Mux_s1_h
    port map (
            O => \N__19441\,
            I => \N__19438\
        );

    \I__4628\ : Span4Mux_h
    port map (
            O => \N__19438\,
            I => \N__19435\
        );

    \I__4627\ : Odrv4
    port map (
            O => \N__19435\,
            I => \GB_BUFFER_SLM_CLK_c_THRU_CO\
        );

    \I__4626\ : InMux
    port map (
            O => \N__19432\,
            I => \N__19429\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__19429\,
            I => \N__19426\
        );

    \I__4624\ : Span4Mux_v
    port map (
            O => \N__19426\,
            I => \N__19423\
        );

    \I__4623\ : IoSpan4Mux
    port map (
            O => \N__19423\,
            I => \N__19420\
        );

    \I__4622\ : Odrv4
    port map (
            O => \N__19420\,
            I => \UART_RX_c\
        );

    \I__4621\ : InMux
    port map (
            O => \N__19417\,
            I => \N__19414\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__19414\,
            I => \N__19411\
        );

    \I__4619\ : Odrv12
    port map (
            O => \N__19411\,
            I => \pc_rx.r_Rx_Data_R\
        );

    \I__4618\ : InMux
    port map (
            O => \N__19408\,
            I => \N__19405\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__19405\,
            I => \N__19395\
        );

    \I__4616\ : ClkMux
    port map (
            O => \N__19404\,
            I => \N__19168\
        );

    \I__4615\ : ClkMux
    port map (
            O => \N__19403\,
            I => \N__19168\
        );

    \I__4614\ : ClkMux
    port map (
            O => \N__19402\,
            I => \N__19168\
        );

    \I__4613\ : ClkMux
    port map (
            O => \N__19401\,
            I => \N__19168\
        );

    \I__4612\ : ClkMux
    port map (
            O => \N__19400\,
            I => \N__19168\
        );

    \I__4611\ : ClkMux
    port map (
            O => \N__19399\,
            I => \N__19168\
        );

    \I__4610\ : ClkMux
    port map (
            O => \N__19398\,
            I => \N__19168\
        );

    \I__4609\ : Glb2LocalMux
    port map (
            O => \N__19395\,
            I => \N__19168\
        );

    \I__4608\ : ClkMux
    port map (
            O => \N__19394\,
            I => \N__19168\
        );

    \I__4607\ : ClkMux
    port map (
            O => \N__19393\,
            I => \N__19168\
        );

    \I__4606\ : ClkMux
    port map (
            O => \N__19392\,
            I => \N__19168\
        );

    \I__4605\ : ClkMux
    port map (
            O => \N__19391\,
            I => \N__19168\
        );

    \I__4604\ : ClkMux
    port map (
            O => \N__19390\,
            I => \N__19168\
        );

    \I__4603\ : ClkMux
    port map (
            O => \N__19389\,
            I => \N__19168\
        );

    \I__4602\ : ClkMux
    port map (
            O => \N__19388\,
            I => \N__19168\
        );

    \I__4601\ : ClkMux
    port map (
            O => \N__19387\,
            I => \N__19168\
        );

    \I__4600\ : ClkMux
    port map (
            O => \N__19386\,
            I => \N__19168\
        );

    \I__4599\ : ClkMux
    port map (
            O => \N__19385\,
            I => \N__19168\
        );

    \I__4598\ : ClkMux
    port map (
            O => \N__19384\,
            I => \N__19168\
        );

    \I__4597\ : ClkMux
    port map (
            O => \N__19383\,
            I => \N__19168\
        );

    \I__4596\ : ClkMux
    port map (
            O => \N__19382\,
            I => \N__19168\
        );

    \I__4595\ : ClkMux
    port map (
            O => \N__19381\,
            I => \N__19168\
        );

    \I__4594\ : ClkMux
    port map (
            O => \N__19380\,
            I => \N__19168\
        );

    \I__4593\ : ClkMux
    port map (
            O => \N__19379\,
            I => \N__19168\
        );

    \I__4592\ : ClkMux
    port map (
            O => \N__19378\,
            I => \N__19168\
        );

    \I__4591\ : ClkMux
    port map (
            O => \N__19377\,
            I => \N__19168\
        );

    \I__4590\ : ClkMux
    port map (
            O => \N__19376\,
            I => \N__19168\
        );

    \I__4589\ : ClkMux
    port map (
            O => \N__19375\,
            I => \N__19168\
        );

    \I__4588\ : ClkMux
    port map (
            O => \N__19374\,
            I => \N__19168\
        );

    \I__4587\ : ClkMux
    port map (
            O => \N__19373\,
            I => \N__19168\
        );

    \I__4586\ : ClkMux
    port map (
            O => \N__19372\,
            I => \N__19168\
        );

    \I__4585\ : ClkMux
    port map (
            O => \N__19371\,
            I => \N__19168\
        );

    \I__4584\ : ClkMux
    port map (
            O => \N__19370\,
            I => \N__19168\
        );

    \I__4583\ : ClkMux
    port map (
            O => \N__19369\,
            I => \N__19168\
        );

    \I__4582\ : ClkMux
    port map (
            O => \N__19368\,
            I => \N__19168\
        );

    \I__4581\ : ClkMux
    port map (
            O => \N__19367\,
            I => \N__19168\
        );

    \I__4580\ : ClkMux
    port map (
            O => \N__19366\,
            I => \N__19168\
        );

    \I__4579\ : ClkMux
    port map (
            O => \N__19365\,
            I => \N__19168\
        );

    \I__4578\ : ClkMux
    port map (
            O => \N__19364\,
            I => \N__19168\
        );

    \I__4577\ : ClkMux
    port map (
            O => \N__19363\,
            I => \N__19168\
        );

    \I__4576\ : ClkMux
    port map (
            O => \N__19362\,
            I => \N__19168\
        );

    \I__4575\ : ClkMux
    port map (
            O => \N__19361\,
            I => \N__19168\
        );

    \I__4574\ : ClkMux
    port map (
            O => \N__19360\,
            I => \N__19168\
        );

    \I__4573\ : ClkMux
    port map (
            O => \N__19359\,
            I => \N__19168\
        );

    \I__4572\ : ClkMux
    port map (
            O => \N__19358\,
            I => \N__19168\
        );

    \I__4571\ : ClkMux
    port map (
            O => \N__19357\,
            I => \N__19168\
        );

    \I__4570\ : ClkMux
    port map (
            O => \N__19356\,
            I => \N__19168\
        );

    \I__4569\ : ClkMux
    port map (
            O => \N__19355\,
            I => \N__19168\
        );

    \I__4568\ : ClkMux
    port map (
            O => \N__19354\,
            I => \N__19168\
        );

    \I__4567\ : ClkMux
    port map (
            O => \N__19353\,
            I => \N__19168\
        );

    \I__4566\ : ClkMux
    port map (
            O => \N__19352\,
            I => \N__19168\
        );

    \I__4565\ : ClkMux
    port map (
            O => \N__19351\,
            I => \N__19168\
        );

    \I__4564\ : ClkMux
    port map (
            O => \N__19350\,
            I => \N__19168\
        );

    \I__4563\ : ClkMux
    port map (
            O => \N__19349\,
            I => \N__19168\
        );

    \I__4562\ : ClkMux
    port map (
            O => \N__19348\,
            I => \N__19168\
        );

    \I__4561\ : ClkMux
    port map (
            O => \N__19347\,
            I => \N__19168\
        );

    \I__4560\ : ClkMux
    port map (
            O => \N__19346\,
            I => \N__19168\
        );

    \I__4559\ : ClkMux
    port map (
            O => \N__19345\,
            I => \N__19168\
        );

    \I__4558\ : ClkMux
    port map (
            O => \N__19344\,
            I => \N__19168\
        );

    \I__4557\ : ClkMux
    port map (
            O => \N__19343\,
            I => \N__19168\
        );

    \I__4556\ : ClkMux
    port map (
            O => \N__19342\,
            I => \N__19168\
        );

    \I__4555\ : ClkMux
    port map (
            O => \N__19341\,
            I => \N__19168\
        );

    \I__4554\ : ClkMux
    port map (
            O => \N__19340\,
            I => \N__19168\
        );

    \I__4553\ : ClkMux
    port map (
            O => \N__19339\,
            I => \N__19168\
        );

    \I__4552\ : ClkMux
    port map (
            O => \N__19338\,
            I => \N__19168\
        );

    \I__4551\ : ClkMux
    port map (
            O => \N__19337\,
            I => \N__19168\
        );

    \I__4550\ : ClkMux
    port map (
            O => \N__19336\,
            I => \N__19168\
        );

    \I__4549\ : ClkMux
    port map (
            O => \N__19335\,
            I => \N__19168\
        );

    \I__4548\ : ClkMux
    port map (
            O => \N__19334\,
            I => \N__19168\
        );

    \I__4547\ : ClkMux
    port map (
            O => \N__19333\,
            I => \N__19168\
        );

    \I__4546\ : ClkMux
    port map (
            O => \N__19332\,
            I => \N__19168\
        );

    \I__4545\ : ClkMux
    port map (
            O => \N__19331\,
            I => \N__19168\
        );

    \I__4544\ : ClkMux
    port map (
            O => \N__19330\,
            I => \N__19168\
        );

    \I__4543\ : ClkMux
    port map (
            O => \N__19329\,
            I => \N__19168\
        );

    \I__4542\ : ClkMux
    port map (
            O => \N__19328\,
            I => \N__19168\
        );

    \I__4541\ : ClkMux
    port map (
            O => \N__19327\,
            I => \N__19168\
        );

    \I__4540\ : ClkMux
    port map (
            O => \N__19326\,
            I => \N__19168\
        );

    \I__4539\ : ClkMux
    port map (
            O => \N__19325\,
            I => \N__19168\
        );

    \I__4538\ : GlobalMux
    port map (
            O => \N__19168\,
            I => \N__19165\
        );

    \I__4537\ : gio2CtrlBuf
    port map (
            O => \N__19165\,
            I => \SLM_CLK_c\
        );

    \I__4536\ : InMux
    port map (
            O => \N__19162\,
            I => \N__19159\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__19159\,
            I => n14
        );

    \I__4534\ : InMux
    port map (
            O => \N__19156\,
            I => n4833
        );

    \I__4533\ : InMux
    port map (
            O => \N__19153\,
            I => \N__19150\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__19150\,
            I => n13
        );

    \I__4531\ : InMux
    port map (
            O => \N__19147\,
            I => n4834
        );

    \I__4530\ : InMux
    port map (
            O => \N__19144\,
            I => \N__19141\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__19141\,
            I => n12
        );

    \I__4528\ : InMux
    port map (
            O => \N__19138\,
            I => n4835
        );

    \I__4527\ : InMux
    port map (
            O => \N__19135\,
            I => \N__19132\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__19132\,
            I => n11_adj_661
        );

    \I__4525\ : InMux
    port map (
            O => \N__19129\,
            I => n4836
        );

    \I__4524\ : InMux
    port map (
            O => \N__19126\,
            I => \N__19123\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__19123\,
            I => n10
        );

    \I__4522\ : InMux
    port map (
            O => \N__19120\,
            I => n4837
        );

    \I__4521\ : InMux
    port map (
            O => \N__19117\,
            I => \N__19114\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__19114\,
            I => n9
        );

    \I__4519\ : InMux
    port map (
            O => \N__19111\,
            I => \bfn_23_7_0_\
        );

    \I__4518\ : InMux
    port map (
            O => \N__19108\,
            I => \N__19105\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__19105\,
            I => n8
        );

    \I__4516\ : InMux
    port map (
            O => \N__19102\,
            I => n4839
        );

    \I__4515\ : InMux
    port map (
            O => \N__19099\,
            I => \N__19096\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__19096\,
            I => n7
        );

    \I__4513\ : InMux
    port map (
            O => \N__19093\,
            I => n4840
        );

    \I__4512\ : InMux
    port map (
            O => \N__19090\,
            I => \N__19087\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__19087\,
            I => n6
        );

    \I__4510\ : InMux
    port map (
            O => \N__19084\,
            I => n4841
        );

    \I__4509\ : InMux
    port map (
            O => \N__19081\,
            I => \N__19078\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__19078\,
            I => n22
        );

    \I__4507\ : InMux
    port map (
            O => \N__19075\,
            I => n4825
        );

    \I__4506\ : InMux
    port map (
            O => \N__19072\,
            I => \N__19069\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__19069\,
            I => n21
        );

    \I__4504\ : InMux
    port map (
            O => \N__19066\,
            I => n4826
        );

    \I__4503\ : InMux
    port map (
            O => \N__19063\,
            I => \N__19060\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__19060\,
            I => n20
        );

    \I__4501\ : InMux
    port map (
            O => \N__19057\,
            I => n4827
        );

    \I__4500\ : InMux
    port map (
            O => \N__19054\,
            I => \N__19051\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__19051\,
            I => n19
        );

    \I__4498\ : InMux
    port map (
            O => \N__19048\,
            I => n4828
        );

    \I__4497\ : InMux
    port map (
            O => \N__19045\,
            I => \N__19042\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__19042\,
            I => n18
        );

    \I__4495\ : InMux
    port map (
            O => \N__19039\,
            I => n4829
        );

    \I__4494\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19033\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__19033\,
            I => n17
        );

    \I__4492\ : InMux
    port map (
            O => \N__19030\,
            I => \bfn_23_6_0_\
        );

    \I__4491\ : InMux
    port map (
            O => \N__19027\,
            I => \N__19024\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__19024\,
            I => n16
        );

    \I__4489\ : InMux
    port map (
            O => \N__19021\,
            I => n4831
        );

    \I__4488\ : InMux
    port map (
            O => \N__19018\,
            I => \N__19015\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__19015\,
            I => n15_adj_663
        );

    \I__4486\ : InMux
    port map (
            O => \N__19012\,
            I => n4832
        );

    \I__4485\ : InMux
    port map (
            O => \N__19009\,
            I => \N__19006\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__19006\,
            I => \N__19003\
        );

    \I__4483\ : Span12Mux_v
    port map (
            O => \N__19003\,
            I => \N__19000\
        );

    \I__4482\ : Span12Mux_v
    port map (
            O => \N__19000\,
            I => \N__18997\
        );

    \I__4481\ : Span12Mux_h
    port map (
            O => \N__18997\,
            I => \N__18994\
        );

    \I__4480\ : Odrv12
    port map (
            O => \N__18994\,
            I => \FIFO_D17_c_17\
        );

    \I__4479\ : IoInMux
    port map (
            O => \N__18991\,
            I => \N__18988\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__18988\,
            I => \N__18985\
        );

    \I__4477\ : Span4Mux_s3_v
    port map (
            O => \N__18985\,
            I => \N__18982\
        );

    \I__4476\ : Span4Mux_v
    port map (
            O => \N__18982\,
            I => \N__18979\
        );

    \I__4475\ : Span4Mux_v
    port map (
            O => \N__18979\,
            I => \N__18976\
        );

    \I__4474\ : Sp12to4
    port map (
            O => \N__18976\,
            I => \N__18973\
        );

    \I__4473\ : Odrv12
    port map (
            O => \N__18973\,
            I => \DATA17_c_17\
        );

    \I__4472\ : InMux
    port map (
            O => \N__18970\,
            I => \N__18966\
        );

    \I__4471\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18963\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__18966\,
            I => \N__18951\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__18963\,
            I => \N__18948\
        );

    \I__4468\ : InMux
    port map (
            O => \N__18962\,
            I => \N__18943\
        );

    \I__4467\ : InMux
    port map (
            O => \N__18961\,
            I => \N__18943\
        );

    \I__4466\ : InMux
    port map (
            O => \N__18960\,
            I => \N__18940\
        );

    \I__4465\ : InMux
    port map (
            O => \N__18959\,
            I => \N__18937\
        );

    \I__4464\ : InMux
    port map (
            O => \N__18958\,
            I => \N__18928\
        );

    \I__4463\ : InMux
    port map (
            O => \N__18957\,
            I => \N__18923\
        );

    \I__4462\ : InMux
    port map (
            O => \N__18956\,
            I => \N__18923\
        );

    \I__4461\ : InMux
    port map (
            O => \N__18955\,
            I => \N__18920\
        );

    \I__4460\ : InMux
    port map (
            O => \N__18954\,
            I => \N__18916\
        );

    \I__4459\ : Span4Mux_v
    port map (
            O => \N__18951\,
            I => \N__18911\
        );

    \I__4458\ : Span4Mux_v
    port map (
            O => \N__18948\,
            I => \N__18904\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__18943\,
            I => \N__18904\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__18940\,
            I => \N__18904\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__18937\,
            I => \N__18901\
        );

    \I__4454\ : InMux
    port map (
            O => \N__18936\,
            I => \N__18898\
        );

    \I__4453\ : InMux
    port map (
            O => \N__18935\,
            I => \N__18893\
        );

    \I__4452\ : InMux
    port map (
            O => \N__18934\,
            I => \N__18893\
        );

    \I__4451\ : InMux
    port map (
            O => \N__18933\,
            I => \N__18890\
        );

    \I__4450\ : InMux
    port map (
            O => \N__18932\,
            I => \N__18887\
        );

    \I__4449\ : InMux
    port map (
            O => \N__18931\,
            I => \N__18883\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__18928\,
            I => \N__18878\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__18923\,
            I => \N__18873\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__18920\,
            I => \N__18873\
        );

    \I__4445\ : InMux
    port map (
            O => \N__18919\,
            I => \N__18867\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__18916\,
            I => \N__18863\
        );

    \I__4443\ : InMux
    port map (
            O => \N__18915\,
            I => \N__18860\
        );

    \I__4442\ : InMux
    port map (
            O => \N__18914\,
            I => \N__18857\
        );

    \I__4441\ : Span4Mux_v
    port map (
            O => \N__18911\,
            I => \N__18852\
        );

    \I__4440\ : Span4Mux_v
    port map (
            O => \N__18904\,
            I => \N__18852\
        );

    \I__4439\ : Span4Mux_h
    port map (
            O => \N__18901\,
            I => \N__18841\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__18898\,
            I => \N__18841\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__18893\,
            I => \N__18841\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__18890\,
            I => \N__18841\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__18887\,
            I => \N__18841\
        );

    \I__4434\ : InMux
    port map (
            O => \N__18886\,
            I => \N__18838\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__18883\,
            I => \N__18835\
        );

    \I__4432\ : InMux
    port map (
            O => \N__18882\,
            I => \N__18832\
        );

    \I__4431\ : InMux
    port map (
            O => \N__18881\,
            I => \N__18829\
        );

    \I__4430\ : Span4Mux_h
    port map (
            O => \N__18878\,
            I => \N__18825\
        );

    \I__4429\ : Span4Mux_v
    port map (
            O => \N__18873\,
            I => \N__18822\
        );

    \I__4428\ : InMux
    port map (
            O => \N__18872\,
            I => \N__18819\
        );

    \I__4427\ : InMux
    port map (
            O => \N__18871\,
            I => \N__18816\
        );

    \I__4426\ : InMux
    port map (
            O => \N__18870\,
            I => \N__18813\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__18867\,
            I => \N__18807\
        );

    \I__4424\ : InMux
    port map (
            O => \N__18866\,
            I => \N__18804\
        );

    \I__4423\ : Span4Mux_v
    port map (
            O => \N__18863\,
            I => \N__18797\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__18860\,
            I => \N__18797\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__18857\,
            I => \N__18797\
        );

    \I__4420\ : Span4Mux_h
    port map (
            O => \N__18852\,
            I => \N__18790\
        );

    \I__4419\ : Span4Mux_v
    port map (
            O => \N__18841\,
            I => \N__18790\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__18838\,
            I => \N__18790\
        );

    \I__4417\ : Span4Mux_v
    port map (
            O => \N__18835\,
            I => \N__18785\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__18832\,
            I => \N__18785\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__18829\,
            I => \N__18782\
        );

    \I__4414\ : InMux
    port map (
            O => \N__18828\,
            I => \N__18779\
        );

    \I__4413\ : Span4Mux_v
    port map (
            O => \N__18825\,
            I => \N__18774\
        );

    \I__4412\ : Span4Mux_h
    port map (
            O => \N__18822\,
            I => \N__18774\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__18819\,
            I => \N__18767\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__18816\,
            I => \N__18767\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__18813\,
            I => \N__18767\
        );

    \I__4408\ : InMux
    port map (
            O => \N__18812\,
            I => \N__18764\
        );

    \I__4407\ : InMux
    port map (
            O => \N__18811\,
            I => \N__18761\
        );

    \I__4406\ : CascadeMux
    port map (
            O => \N__18810\,
            I => \N__18755\
        );

    \I__4405\ : Span4Mux_v
    port map (
            O => \N__18807\,
            I => \N__18752\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__18804\,
            I => \N__18749\
        );

    \I__4403\ : Span4Mux_v
    port map (
            O => \N__18797\,
            I => \N__18742\
        );

    \I__4402\ : Span4Mux_h
    port map (
            O => \N__18790\,
            I => \N__18742\
        );

    \I__4401\ : Span4Mux_v
    port map (
            O => \N__18785\,
            I => \N__18742\
        );

    \I__4400\ : Span12Mux_h
    port map (
            O => \N__18782\,
            I => \N__18737\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__18779\,
            I => \N__18737\
        );

    \I__4398\ : Span4Mux_h
    port map (
            O => \N__18774\,
            I => \N__18728\
        );

    \I__4397\ : Span4Mux_v
    port map (
            O => \N__18767\,
            I => \N__18728\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__18764\,
            I => \N__18728\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__18761\,
            I => \N__18728\
        );

    \I__4394\ : InMux
    port map (
            O => \N__18760\,
            I => \N__18723\
        );

    \I__4393\ : InMux
    port map (
            O => \N__18759\,
            I => \N__18723\
        );

    \I__4392\ : InMux
    port map (
            O => \N__18758\,
            I => \N__18720\
        );

    \I__4391\ : InMux
    port map (
            O => \N__18755\,
            I => \N__18717\
        );

    \I__4390\ : Odrv4
    port map (
            O => \N__18752\,
            I => \bluejay_data_inst.data_output_active_cmd\
        );

    \I__4389\ : Odrv4
    port map (
            O => \N__18749\,
            I => \bluejay_data_inst.data_output_active_cmd\
        );

    \I__4388\ : Odrv4
    port map (
            O => \N__18742\,
            I => \bluejay_data_inst.data_output_active_cmd\
        );

    \I__4387\ : Odrv12
    port map (
            O => \N__18737\,
            I => \bluejay_data_inst.data_output_active_cmd\
        );

    \I__4386\ : Odrv4
    port map (
            O => \N__18728\,
            I => \bluejay_data_inst.data_output_active_cmd\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__18723\,
            I => \bluejay_data_inst.data_output_active_cmd\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__18720\,
            I => \bluejay_data_inst.data_output_active_cmd\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__18717\,
            I => \bluejay_data_inst.data_output_active_cmd\
        );

    \I__4382\ : InMux
    port map (
            O => \N__18700\,
            I => \N__18697\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__18697\,
            I => \N__18694\
        );

    \I__4380\ : Span4Mux_v
    port map (
            O => \N__18694\,
            I => \N__18691\
        );

    \I__4379\ : Sp12to4
    port map (
            O => \N__18691\,
            I => \N__18688\
        );

    \I__4378\ : Span12Mux_s8_h
    port map (
            O => \N__18688\,
            I => \N__18685\
        );

    \I__4377\ : Span12Mux_v
    port map (
            O => \N__18685\,
            I => \N__18682\
        );

    \I__4376\ : Odrv12
    port map (
            O => \N__18682\,
            I => \FIFO_D2_c_2\
        );

    \I__4375\ : IoInMux
    port map (
            O => \N__18679\,
            I => \N__18676\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__18676\,
            I => \N__18673\
        );

    \I__4373\ : Span12Mux_s10_v
    port map (
            O => \N__18673\,
            I => \N__18670\
        );

    \I__4372\ : Odrv12
    port map (
            O => \N__18670\,
            I => \DATA2_c_2\
        );

    \I__4371\ : InMux
    port map (
            O => \N__18667\,
            I => \N__18664\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__18664\,
            I => \N__18660\
        );

    \I__4369\ : InMux
    port map (
            O => \N__18663\,
            I => \N__18657\
        );

    \I__4368\ : Span12Mux_s7_h
    port map (
            O => \N__18660\,
            I => \N__18652\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__18657\,
            I => \N__18649\
        );

    \I__4366\ : InMux
    port map (
            O => \N__18656\,
            I => \N__18646\
        );

    \I__4365\ : InMux
    port map (
            O => \N__18655\,
            I => \N__18643\
        );

    \I__4364\ : Span12Mux_h
    port map (
            O => \N__18652\,
            I => \N__18640\
        );

    \I__4363\ : Span4Mux_v
    port map (
            O => \N__18649\,
            I => \N__18637\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__18646\,
            I => \N__18634\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__18643\,
            I => \N__18631\
        );

    \I__4360\ : Odrv12
    port map (
            O => \N__18640\,
            I => get_next_word_cmd
        );

    \I__4359\ : Odrv4
    port map (
            O => \N__18637\,
            I => get_next_word_cmd
        );

    \I__4358\ : Odrv4
    port map (
            O => \N__18634\,
            I => get_next_word_cmd
        );

    \I__4357\ : Odrv4
    port map (
            O => \N__18631\,
            I => get_next_word_cmd
        );

    \I__4356\ : IoInMux
    port map (
            O => \N__18622\,
            I => \N__18619\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__18619\,
            I => \N__18616\
        );

    \I__4354\ : Span4Mux_s2_v
    port map (
            O => \N__18616\,
            I => \N__18613\
        );

    \I__4353\ : Sp12to4
    port map (
            O => \N__18613\,
            I => \N__18610\
        );

    \I__4352\ : Span12Mux_s9_h
    port map (
            O => \N__18610\,
            I => \N__18607\
        );

    \I__4351\ : Odrv12
    port map (
            O => \N__18607\,
            I => \DEBUG_8_c\
        );

    \I__4350\ : InMux
    port map (
            O => \N__18604\,
            I => \N__18597\
        );

    \I__4349\ : InMux
    port map (
            O => \N__18603\,
            I => \N__18588\
        );

    \I__4348\ : InMux
    port map (
            O => \N__18602\,
            I => \N__18584\
        );

    \I__4347\ : InMux
    port map (
            O => \N__18601\,
            I => \N__18581\
        );

    \I__4346\ : InMux
    port map (
            O => \N__18600\,
            I => \N__18572\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__18597\,
            I => \N__18569\
        );

    \I__4344\ : InMux
    port map (
            O => \N__18596\,
            I => \N__18564\
        );

    \I__4343\ : InMux
    port map (
            O => \N__18595\,
            I => \N__18564\
        );

    \I__4342\ : InMux
    port map (
            O => \N__18594\,
            I => \N__18559\
        );

    \I__4341\ : InMux
    port map (
            O => \N__18593\,
            I => \N__18559\
        );

    \I__4340\ : InMux
    port map (
            O => \N__18592\,
            I => \N__18556\
        );

    \I__4339\ : InMux
    port map (
            O => \N__18591\,
            I => \N__18553\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__18588\,
            I => \N__18550\
        );

    \I__4337\ : InMux
    port map (
            O => \N__18587\,
            I => \N__18547\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__18584\,
            I => \N__18539\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__18581\,
            I => \N__18539\
        );

    \I__4334\ : InMux
    port map (
            O => \N__18580\,
            I => \N__18536\
        );

    \I__4333\ : InMux
    port map (
            O => \N__18579\,
            I => \N__18525\
        );

    \I__4332\ : InMux
    port map (
            O => \N__18578\,
            I => \N__18525\
        );

    \I__4331\ : InMux
    port map (
            O => \N__18577\,
            I => \N__18525\
        );

    \I__4330\ : InMux
    port map (
            O => \N__18576\,
            I => \N__18525\
        );

    \I__4329\ : InMux
    port map (
            O => \N__18575\,
            I => \N__18525\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__18572\,
            I => \N__18522\
        );

    \I__4327\ : Span4Mux_h
    port map (
            O => \N__18569\,
            I => \N__18515\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__18564\,
            I => \N__18515\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__18559\,
            I => \N__18515\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__18556\,
            I => \N__18510\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__18553\,
            I => \N__18510\
        );

    \I__4322\ : Span4Mux_h
    port map (
            O => \N__18550\,
            I => \N__18501\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__18547\,
            I => \N__18498\
        );

    \I__4320\ : InMux
    port map (
            O => \N__18546\,
            I => \N__18495\
        );

    \I__4319\ : InMux
    port map (
            O => \N__18545\,
            I => \N__18490\
        );

    \I__4318\ : InMux
    port map (
            O => \N__18544\,
            I => \N__18490\
        );

    \I__4317\ : Span4Mux_h
    port map (
            O => \N__18539\,
            I => \N__18487\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__18536\,
            I => \N__18482\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__18525\,
            I => \N__18482\
        );

    \I__4314\ : Span4Mux_h
    port map (
            O => \N__18522\,
            I => \N__18475\
        );

    \I__4313\ : Span4Mux_h
    port map (
            O => \N__18515\,
            I => \N__18475\
        );

    \I__4312\ : Span4Mux_h
    port map (
            O => \N__18510\,
            I => \N__18475\
        );

    \I__4311\ : InMux
    port map (
            O => \N__18509\,
            I => \N__18472\
        );

    \I__4310\ : InMux
    port map (
            O => \N__18508\,
            I => \N__18467\
        );

    \I__4309\ : InMux
    port map (
            O => \N__18507\,
            I => \N__18467\
        );

    \I__4308\ : InMux
    port map (
            O => \N__18506\,
            I => \N__18462\
        );

    \I__4307\ : InMux
    port map (
            O => \N__18505\,
            I => \N__18462\
        );

    \I__4306\ : InMux
    port map (
            O => \N__18504\,
            I => \N__18459\
        );

    \I__4305\ : Odrv4
    port map (
            O => \N__18501\,
            I => state_2
        );

    \I__4304\ : Odrv4
    port map (
            O => \N__18498\,
            I => state_2
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__18495\,
            I => state_2
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__18490\,
            I => state_2
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__18487\,
            I => state_2
        );

    \I__4300\ : Odrv12
    port map (
            O => \N__18482\,
            I => state_2
        );

    \I__4299\ : Odrv4
    port map (
            O => \N__18475\,
            I => state_2
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__18472\,
            I => state_2
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__18467\,
            I => state_2
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__18462\,
            I => state_2
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__18459\,
            I => state_2
        );

    \I__4294\ : InMux
    port map (
            O => \N__18436\,
            I => \N__18420\
        );

    \I__4293\ : CascadeMux
    port map (
            O => \N__18435\,
            I => \N__18415\
        );

    \I__4292\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18410\
        );

    \I__4291\ : InMux
    port map (
            O => \N__18433\,
            I => \N__18407\
        );

    \I__4290\ : InMux
    port map (
            O => \N__18432\,
            I => \N__18404\
        );

    \I__4289\ : InMux
    port map (
            O => \N__18431\,
            I => \N__18401\
        );

    \I__4288\ : InMux
    port map (
            O => \N__18430\,
            I => \N__18396\
        );

    \I__4287\ : InMux
    port map (
            O => \N__18429\,
            I => \N__18396\
        );

    \I__4286\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18391\
        );

    \I__4285\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18391\
        );

    \I__4284\ : InMux
    port map (
            O => \N__18426\,
            I => \N__18381\
        );

    \I__4283\ : InMux
    port map (
            O => \N__18425\,
            I => \N__18381\
        );

    \I__4282\ : InMux
    port map (
            O => \N__18424\,
            I => \N__18381\
        );

    \I__4281\ : InMux
    port map (
            O => \N__18423\,
            I => \N__18376\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__18420\,
            I => \N__18373\
        );

    \I__4279\ : InMux
    port map (
            O => \N__18419\,
            I => \N__18366\
        );

    \I__4278\ : InMux
    port map (
            O => \N__18418\,
            I => \N__18366\
        );

    \I__4277\ : InMux
    port map (
            O => \N__18415\,
            I => \N__18361\
        );

    \I__4276\ : InMux
    port map (
            O => \N__18414\,
            I => \N__18358\
        );

    \I__4275\ : InMux
    port map (
            O => \N__18413\,
            I => \N__18355\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__18410\,
            I => \N__18352\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__18407\,
            I => \N__18349\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__18404\,
            I => \N__18340\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__18401\,
            I => \N__18340\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__18396\,
            I => \N__18340\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__18391\,
            I => \N__18340\
        );

    \I__4268\ : InMux
    port map (
            O => \N__18390\,
            I => \N__18335\
        );

    \I__4267\ : InMux
    port map (
            O => \N__18389\,
            I => \N__18335\
        );

    \I__4266\ : InMux
    port map (
            O => \N__18388\,
            I => \N__18332\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__18381\,
            I => \N__18329\
        );

    \I__4264\ : InMux
    port map (
            O => \N__18380\,
            I => \N__18324\
        );

    \I__4263\ : InMux
    port map (
            O => \N__18379\,
            I => \N__18324\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__18376\,
            I => \N__18321\
        );

    \I__4261\ : Span4Mux_v
    port map (
            O => \N__18373\,
            I => \N__18318\
        );

    \I__4260\ : InMux
    port map (
            O => \N__18372\,
            I => \N__18315\
        );

    \I__4259\ : InMux
    port map (
            O => \N__18371\,
            I => \N__18312\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__18366\,
            I => \N__18309\
        );

    \I__4257\ : InMux
    port map (
            O => \N__18365\,
            I => \N__18304\
        );

    \I__4256\ : InMux
    port map (
            O => \N__18364\,
            I => \N__18304\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__18361\,
            I => \N__18285\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__18358\,
            I => \N__18285\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__18355\,
            I => \N__18285\
        );

    \I__4252\ : Span4Mux_v
    port map (
            O => \N__18352\,
            I => \N__18285\
        );

    \I__4251\ : Span4Mux_v
    port map (
            O => \N__18349\,
            I => \N__18285\
        );

    \I__4250\ : Span4Mux_v
    port map (
            O => \N__18340\,
            I => \N__18285\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__18335\,
            I => \N__18285\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__18332\,
            I => \N__18285\
        );

    \I__4247\ : Span4Mux_v
    port map (
            O => \N__18329\,
            I => \N__18285\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__18324\,
            I => \bluejay_data_inst.state_1\
        );

    \I__4245\ : Odrv4
    port map (
            O => \N__18321\,
            I => \bluejay_data_inst.state_1\
        );

    \I__4244\ : Odrv4
    port map (
            O => \N__18318\,
            I => \bluejay_data_inst.state_1\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__18315\,
            I => \bluejay_data_inst.state_1\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__18312\,
            I => \bluejay_data_inst.state_1\
        );

    \I__4241\ : Odrv4
    port map (
            O => \N__18309\,
            I => \bluejay_data_inst.state_1\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__18304\,
            I => \bluejay_data_inst.state_1\
        );

    \I__4239\ : Odrv4
    port map (
            O => \N__18285\,
            I => \bluejay_data_inst.state_1\
        );

    \I__4238\ : InMux
    port map (
            O => \N__18268\,
            I => \N__18259\
        );

    \I__4237\ : CascadeMux
    port map (
            O => \N__18267\,
            I => \N__18252\
        );

    \I__4236\ : CascadeMux
    port map (
            O => \N__18266\,
            I => \N__18249\
        );

    \I__4235\ : CascadeMux
    port map (
            O => \N__18265\,
            I => \N__18246\
        );

    \I__4234\ : InMux
    port map (
            O => \N__18264\,
            I => \N__18239\
        );

    \I__4233\ : InMux
    port map (
            O => \N__18263\,
            I => \N__18234\
        );

    \I__4232\ : InMux
    port map (
            O => \N__18262\,
            I => \N__18234\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__18259\,
            I => \N__18228\
        );

    \I__4230\ : InMux
    port map (
            O => \N__18258\,
            I => \N__18225\
        );

    \I__4229\ : InMux
    port map (
            O => \N__18257\,
            I => \N__18220\
        );

    \I__4228\ : InMux
    port map (
            O => \N__18256\,
            I => \N__18220\
        );

    \I__4227\ : InMux
    port map (
            O => \N__18255\,
            I => \N__18213\
        );

    \I__4226\ : InMux
    port map (
            O => \N__18252\,
            I => \N__18213\
        );

    \I__4225\ : InMux
    port map (
            O => \N__18249\,
            I => \N__18213\
        );

    \I__4224\ : InMux
    port map (
            O => \N__18246\,
            I => \N__18210\
        );

    \I__4223\ : InMux
    port map (
            O => \N__18245\,
            I => \N__18207\
        );

    \I__4222\ : InMux
    port map (
            O => \N__18244\,
            I => \N__18201\
        );

    \I__4221\ : InMux
    port map (
            O => \N__18243\,
            I => \N__18195\
        );

    \I__4220\ : InMux
    port map (
            O => \N__18242\,
            I => \N__18195\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__18239\,
            I => \N__18192\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__18234\,
            I => \N__18189\
        );

    \I__4217\ : InMux
    port map (
            O => \N__18233\,
            I => \N__18182\
        );

    \I__4216\ : InMux
    port map (
            O => \N__18232\,
            I => \N__18182\
        );

    \I__4215\ : InMux
    port map (
            O => \N__18231\,
            I => \N__18182\
        );

    \I__4214\ : Span4Mux_h
    port map (
            O => \N__18228\,
            I => \N__18172\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__18225\,
            I => \N__18172\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__18220\,
            I => \N__18172\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__18213\,
            I => \N__18169\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__18210\,
            I => \N__18162\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__18207\,
            I => \N__18162\
        );

    \I__4208\ : InMux
    port map (
            O => \N__18206\,
            I => \N__18155\
        );

    \I__4207\ : InMux
    port map (
            O => \N__18205\,
            I => \N__18155\
        );

    \I__4206\ : InMux
    port map (
            O => \N__18204\,
            I => \N__18155\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__18201\,
            I => \N__18152\
        );

    \I__4204\ : InMux
    port map (
            O => \N__18200\,
            I => \N__18149\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__18195\,
            I => \N__18140\
        );

    \I__4202\ : Span4Mux_h
    port map (
            O => \N__18192\,
            I => \N__18140\
        );

    \I__4201\ : Span4Mux_v
    port map (
            O => \N__18189\,
            I => \N__18140\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__18182\,
            I => \N__18140\
        );

    \I__4199\ : InMux
    port map (
            O => \N__18181\,
            I => \N__18137\
        );

    \I__4198\ : InMux
    port map (
            O => \N__18180\,
            I => \N__18132\
        );

    \I__4197\ : InMux
    port map (
            O => \N__18179\,
            I => \N__18132\
        );

    \I__4196\ : Span4Mux_h
    port map (
            O => \N__18172\,
            I => \N__18127\
        );

    \I__4195\ : Span4Mux_h
    port map (
            O => \N__18169\,
            I => \N__18127\
        );

    \I__4194\ : InMux
    port map (
            O => \N__18168\,
            I => \N__18122\
        );

    \I__4193\ : InMux
    port map (
            O => \N__18167\,
            I => \N__18122\
        );

    \I__4192\ : Odrv4
    port map (
            O => \N__18162\,
            I => state_0
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__18155\,
            I => state_0
        );

    \I__4190\ : Odrv4
    port map (
            O => \N__18152\,
            I => state_0
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__18149\,
            I => state_0
        );

    \I__4188\ : Odrv4
    port map (
            O => \N__18140\,
            I => state_0
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__18137\,
            I => state_0
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__18132\,
            I => state_0
        );

    \I__4185\ : Odrv4
    port map (
            O => \N__18127\,
            I => state_0
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__18122\,
            I => state_0
        );

    \I__4183\ : IoInMux
    port map (
            O => \N__18103\,
            I => \N__18100\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__18100\,
            I => \N__18097\
        );

    \I__4181\ : Span12Mux_s4_h
    port map (
            O => \N__18097\,
            I => \N__18094\
        );

    \I__4180\ : Odrv12
    port map (
            O => \N__18094\,
            I => \UPDATE_c\
        );

    \I__4179\ : SRMux
    port map (
            O => \N__18091\,
            I => \N__18088\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__18088\,
            I => \N__18085\
        );

    \I__4177\ : Span4Mux_h
    port map (
            O => \N__18085\,
            I => \N__18082\
        );

    \I__4176\ : Odrv4
    port map (
            O => \N__18082\,
            I => \bluejay_data_inst.n2096\
        );

    \I__4175\ : InMux
    port map (
            O => \N__18079\,
            I => \N__18076\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__18076\,
            I => \N__18068\
        );

    \I__4173\ : InMux
    port map (
            O => \N__18075\,
            I => \N__18065\
        );

    \I__4172\ : InMux
    port map (
            O => \N__18074\,
            I => \N__18060\
        );

    \I__4171\ : InMux
    port map (
            O => \N__18073\,
            I => \N__18060\
        );

    \I__4170\ : InMux
    port map (
            O => \N__18072\,
            I => \N__18055\
        );

    \I__4169\ : InMux
    port map (
            O => \N__18071\,
            I => \N__18055\
        );

    \I__4168\ : Span4Mux_v
    port map (
            O => \N__18068\,
            I => \N__18050\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__18065\,
            I => \N__18047\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__18060\,
            I => \N__18042\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__18055\,
            I => \N__18042\
        );

    \I__4164\ : InMux
    port map (
            O => \N__18054\,
            I => \N__18033\
        );

    \I__4163\ : InMux
    port map (
            O => \N__18053\,
            I => \N__18033\
        );

    \I__4162\ : Span4Mux_h
    port map (
            O => \N__18050\,
            I => \N__18028\
        );

    \I__4161\ : Span4Mux_v
    port map (
            O => \N__18047\,
            I => \N__18028\
        );

    \I__4160\ : Span4Mux_v
    port map (
            O => \N__18042\,
            I => \N__18025\
        );

    \I__4159\ : InMux
    port map (
            O => \N__18041\,
            I => \N__18020\
        );

    \I__4158\ : InMux
    port map (
            O => \N__18040\,
            I => \N__18020\
        );

    \I__4157\ : InMux
    port map (
            O => \N__18039\,
            I => \N__18015\
        );

    \I__4156\ : InMux
    port map (
            O => \N__18038\,
            I => \N__18015\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__18033\,
            I => \N__18012\
        );

    \I__4154\ : Sp12to4
    port map (
            O => \N__18028\,
            I => \N__18001\
        );

    \I__4153\ : Sp12to4
    port map (
            O => \N__18025\,
            I => \N__18001\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__18020\,
            I => \N__18001\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__18015\,
            I => \N__18001\
        );

    \I__4150\ : Span12Mux_v
    port map (
            O => \N__18012\,
            I => \N__18001\
        );

    \I__4149\ : Odrv12
    port map (
            O => \N__18001\,
            I => \r_Rx_Data\
        );

    \I__4148\ : InMux
    port map (
            O => \N__17998\,
            I => \N__17995\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__17995\,
            I => n25_adj_662
        );

    \I__4146\ : InMux
    port map (
            O => \N__17992\,
            I => \bfn_23_5_0_\
        );

    \I__4145\ : InMux
    port map (
            O => \N__17989\,
            I => \N__17986\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__17986\,
            I => n24
        );

    \I__4143\ : InMux
    port map (
            O => \N__17983\,
            I => n4823
        );

    \I__4142\ : InMux
    port map (
            O => \N__17980\,
            I => \N__17977\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__17977\,
            I => n23
        );

    \I__4140\ : InMux
    port map (
            O => \N__17974\,
            I => n4824
        );

    \I__4139\ : CascadeMux
    port map (
            O => \N__17971\,
            I => \N__17964\
        );

    \I__4138\ : InMux
    port map (
            O => \N__17970\,
            I => \N__17961\
        );

    \I__4137\ : InMux
    port map (
            O => \N__17969\,
            I => \N__17956\
        );

    \I__4136\ : InMux
    port map (
            O => \N__17968\,
            I => \N__17956\
        );

    \I__4135\ : InMux
    port map (
            O => \N__17967\,
            I => \N__17953\
        );

    \I__4134\ : InMux
    port map (
            O => \N__17964\,
            I => \N__17950\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__17961\,
            I => \bluejay_data_inst.state_timeout_counter_6\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__17956\,
            I => \bluejay_data_inst.state_timeout_counter_6\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__17953\,
            I => \bluejay_data_inst.state_timeout_counter_6\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__17950\,
            I => \bluejay_data_inst.state_timeout_counter_6\
        );

    \I__4129\ : CascadeMux
    port map (
            O => \N__17941\,
            I => \bluejay_data_inst.state_timeout_counter_7_N_122_6_cascade_\
        );

    \I__4128\ : InMux
    port map (
            O => \N__17938\,
            I => \N__17935\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__17935\,
            I => \bluejay_data_inst.state_timeout_counter_7_N_122_6\
        );

    \I__4126\ : CascadeMux
    port map (
            O => \N__17932\,
            I => \bluejay_data_inst.n8_adj_638_cascade_\
        );

    \I__4125\ : SRMux
    port map (
            O => \N__17929\,
            I => \N__17926\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__17926\,
            I => \N__17923\
        );

    \I__4123\ : Span4Mux_h
    port map (
            O => \N__17923\,
            I => \N__17920\
        );

    \I__4122\ : Odrv4
    port map (
            O => \N__17920\,
            I => \bluejay_data_inst.n4_adj_639\
        );

    \I__4121\ : InMux
    port map (
            O => \N__17917\,
            I => \N__17911\
        );

    \I__4120\ : InMux
    port map (
            O => \N__17916\,
            I => \N__17911\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__17911\,
            I => \N__17908\
        );

    \I__4118\ : Span4Mux_v
    port map (
            O => \N__17908\,
            I => \N__17896\
        );

    \I__4117\ : InMux
    port map (
            O => \N__17907\,
            I => \N__17891\
        );

    \I__4116\ : InMux
    port map (
            O => \N__17906\,
            I => \N__17891\
        );

    \I__4115\ : InMux
    port map (
            O => \N__17905\,
            I => \N__17888\
        );

    \I__4114\ : InMux
    port map (
            O => \N__17904\,
            I => \N__17885\
        );

    \I__4113\ : InMux
    port map (
            O => \N__17903\,
            I => \N__17882\
        );

    \I__4112\ : InMux
    port map (
            O => \N__17902\,
            I => \N__17875\
        );

    \I__4111\ : InMux
    port map (
            O => \N__17901\,
            I => \N__17875\
        );

    \I__4110\ : InMux
    port map (
            O => \N__17900\,
            I => \N__17875\
        );

    \I__4109\ : InMux
    port map (
            O => \N__17899\,
            I => \N__17872\
        );

    \I__4108\ : Sp12to4
    port map (
            O => \N__17896\,
            I => \N__17869\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__17891\,
            I => \N__17866\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__17888\,
            I => \N__17857\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__17885\,
            I => \N__17857\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__17882\,
            I => \N__17857\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__17875\,
            I => \N__17857\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__17872\,
            I => \bluejay_data_inst.n1054\
        );

    \I__4101\ : Odrv12
    port map (
            O => \N__17869\,
            I => \bluejay_data_inst.n1054\
        );

    \I__4100\ : Odrv4
    port map (
            O => \N__17866\,
            I => \bluejay_data_inst.n1054\
        );

    \I__4099\ : Odrv4
    port map (
            O => \N__17857\,
            I => \bluejay_data_inst.n1054\
        );

    \I__4098\ : InMux
    port map (
            O => \N__17848\,
            I => \N__17845\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__17845\,
            I => \bluejay_data_inst.n5521\
        );

    \I__4096\ : InMux
    port map (
            O => \N__17842\,
            I => \N__17838\
        );

    \I__4095\ : InMux
    port map (
            O => \N__17841\,
            I => \N__17833\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__17838\,
            I => \N__17830\
        );

    \I__4093\ : InMux
    port map (
            O => \N__17837\,
            I => \N__17827\
        );

    \I__4092\ : InMux
    port map (
            O => \N__17836\,
            I => \N__17824\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__17833\,
            I => \N__17820\
        );

    \I__4090\ : Span4Mux_h
    port map (
            O => \N__17830\,
            I => \N__17813\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__17827\,
            I => \N__17813\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__17824\,
            I => \N__17813\
        );

    \I__4087\ : InMux
    port map (
            O => \N__17823\,
            I => \N__17810\
        );

    \I__4086\ : Odrv4
    port map (
            O => \N__17820\,
            I => \bluejay_data_inst.n34\
        );

    \I__4085\ : Odrv4
    port map (
            O => \N__17813\,
            I => \bluejay_data_inst.n34\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__17810\,
            I => \bluejay_data_inst.n34\
        );

    \I__4083\ : CascadeMux
    port map (
            O => \N__17803\,
            I => \bluejay_data_inst.state_timeout_counter_7_N_122_0_cascade_\
        );

    \I__4082\ : CascadeMux
    port map (
            O => \N__17800\,
            I => \bluejay_data_inst.n8_adj_645_cascade_\
        );

    \I__4081\ : InMux
    port map (
            O => \N__17797\,
            I => \N__17794\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__17794\,
            I => \bluejay_data_inst.state_timeout_counter_7_N_122_0\
        );

    \I__4079\ : InMux
    port map (
            O => \N__17791\,
            I => \N__17788\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__17788\,
            I => \N__17785\
        );

    \I__4077\ : Odrv12
    port map (
            O => \N__17785\,
            I => \bluejay_data_inst.state_timeout_counter_7_N_122_2\
        );

    \I__4076\ : CascadeMux
    port map (
            O => \N__17782\,
            I => \N__17777\
        );

    \I__4075\ : CascadeMux
    port map (
            O => \N__17781\,
            I => \N__17774\
        );

    \I__4074\ : InMux
    port map (
            O => \N__17780\,
            I => \N__17767\
        );

    \I__4073\ : InMux
    port map (
            O => \N__17777\,
            I => \N__17767\
        );

    \I__4072\ : InMux
    port map (
            O => \N__17774\,
            I => \N__17764\
        );

    \I__4071\ : CascadeMux
    port map (
            O => \N__17773\,
            I => \N__17761\
        );

    \I__4070\ : InMux
    port map (
            O => \N__17772\,
            I => \N__17758\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__17767\,
            I => \N__17755\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__17764\,
            I => \N__17752\
        );

    \I__4067\ : InMux
    port map (
            O => \N__17761\,
            I => \N__17749\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__17758\,
            I => \N__17746\
        );

    \I__4065\ : Span4Mux_v
    port map (
            O => \N__17755\,
            I => \N__17741\
        );

    \I__4064\ : Span4Mux_h
    port map (
            O => \N__17752\,
            I => \N__17741\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__17749\,
            I => n3_adj_669
        );

    \I__4062\ : Odrv4
    port map (
            O => \N__17746\,
            I => n3_adj_669
        );

    \I__4061\ : Odrv4
    port map (
            O => \N__17741\,
            I => n3_adj_669
        );

    \I__4060\ : InMux
    port map (
            O => \N__17734\,
            I => \N__17731\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__17731\,
            I => \N__17728\
        );

    \I__4058\ : Odrv12
    port map (
            O => \N__17728\,
            I => \bluejay_data_inst.n4260\
        );

    \I__4057\ : InMux
    port map (
            O => \N__17725\,
            I => \N__17722\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__17722\,
            I => \N__17718\
        );

    \I__4055\ : InMux
    port map (
            O => \N__17721\,
            I => \N__17715\
        );

    \I__4054\ : Span4Mux_v
    port map (
            O => \N__17718\,
            I => \N__17708\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__17715\,
            I => \N__17708\
        );

    \I__4052\ : InMux
    port map (
            O => \N__17714\,
            I => \N__17705\
        );

    \I__4051\ : InMux
    port map (
            O => \N__17713\,
            I => \N__17701\
        );

    \I__4050\ : Span4Mux_h
    port map (
            O => \N__17708\,
            I => \N__17698\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__17705\,
            I => \N__17695\
        );

    \I__4048\ : InMux
    port map (
            O => \N__17704\,
            I => \N__17692\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__17701\,
            I => \bluejay_data_inst.state_timeout_counter_2\
        );

    \I__4046\ : Odrv4
    port map (
            O => \N__17698\,
            I => \bluejay_data_inst.state_timeout_counter_2\
        );

    \I__4045\ : Odrv4
    port map (
            O => \N__17695\,
            I => \bluejay_data_inst.state_timeout_counter_2\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__17692\,
            I => \bluejay_data_inst.state_timeout_counter_2\
        );

    \I__4043\ : SRMux
    port map (
            O => \N__17683\,
            I => \N__17680\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__17680\,
            I => \N__17677\
        );

    \I__4041\ : Odrv12
    port map (
            O => \N__17677\,
            I => \bluejay_data_inst.n4_adj_650\
        );

    \I__4040\ : InMux
    port map (
            O => \N__17674\,
            I => \N__17666\
        );

    \I__4039\ : InMux
    port map (
            O => \N__17673\,
            I => \N__17666\
        );

    \I__4038\ : InMux
    port map (
            O => \N__17672\,
            I => \N__17663\
        );

    \I__4037\ : InMux
    port map (
            O => \N__17671\,
            I => \N__17660\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__17666\,
            I => \N__17652\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__17663\,
            I => \N__17652\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__17660\,
            I => \N__17652\
        );

    \I__4033\ : InMux
    port map (
            O => \N__17659\,
            I => \N__17649\
        );

    \I__4032\ : Span4Mux_v
    port map (
            O => \N__17652\,
            I => \N__17646\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__17649\,
            I => \bluejay_data_inst.state_timeout_counter_0\
        );

    \I__4030\ : Odrv4
    port map (
            O => \N__17646\,
            I => \bluejay_data_inst.state_timeout_counter_0\
        );

    \I__4029\ : SRMux
    port map (
            O => \N__17641\,
            I => \N__17638\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__17638\,
            I => \N__17635\
        );

    \I__4027\ : Span4Mux_v
    port map (
            O => \N__17635\,
            I => \N__17632\
        );

    \I__4026\ : Odrv4
    port map (
            O => \N__17632\,
            I => \bluejay_data_inst.n4_adj_636\
        );

    \I__4025\ : InMux
    port map (
            O => \N__17629\,
            I => \N__17626\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__17626\,
            I => \N__17623\
        );

    \I__4023\ : Span4Mux_v
    port map (
            O => \N__17623\,
            I => \N__17620\
        );

    \I__4022\ : Sp12to4
    port map (
            O => \N__17620\,
            I => \N__17617\
        );

    \I__4021\ : Span12Mux_h
    port map (
            O => \N__17617\,
            I => \N__17614\
        );

    \I__4020\ : Span12Mux_v
    port map (
            O => \N__17614\,
            I => \N__17611\
        );

    \I__4019\ : Odrv12
    port map (
            O => \N__17611\,
            I => \FIFO_D7_c_7\
        );

    \I__4018\ : IoInMux
    port map (
            O => \N__17608\,
            I => \N__17605\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__17605\,
            I => \N__17602\
        );

    \I__4016\ : Span4Mux_s3_h
    port map (
            O => \N__17602\,
            I => \N__17599\
        );

    \I__4015\ : Span4Mux_h
    port map (
            O => \N__17599\,
            I => \N__17596\
        );

    \I__4014\ : Sp12to4
    port map (
            O => \N__17596\,
            I => \N__17593\
        );

    \I__4013\ : Span12Mux_v
    port map (
            O => \N__17593\,
            I => \N__17590\
        );

    \I__4012\ : Odrv12
    port map (
            O => \N__17590\,
            I => \DATA7_c_7\
        );

    \I__4011\ : InMux
    port map (
            O => \N__17587\,
            I => \N__17581\
        );

    \I__4010\ : InMux
    port map (
            O => \N__17586\,
            I => \N__17573\
        );

    \I__4009\ : InMux
    port map (
            O => \N__17585\,
            I => \N__17573\
        );

    \I__4008\ : InMux
    port map (
            O => \N__17584\,
            I => \N__17573\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__17581\,
            I => \N__17570\
        );

    \I__4006\ : InMux
    port map (
            O => \N__17580\,
            I => \N__17567\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__17573\,
            I => \bluejay_data_inst.state_timeout_counter_7\
        );

    \I__4004\ : Odrv4
    port map (
            O => \N__17570\,
            I => \bluejay_data_inst.state_timeout_counter_7\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__17567\,
            I => \bluejay_data_inst.state_timeout_counter_7\
        );

    \I__4002\ : SRMux
    port map (
            O => \N__17560\,
            I => \N__17557\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__17557\,
            I => \N__17554\
        );

    \I__4000\ : Odrv4
    port map (
            O => \N__17554\,
            I => \bluejay_data_inst.n4_adj_641\
        );

    \I__3999\ : InMux
    port map (
            O => \N__17551\,
            I => \N__17544\
        );

    \I__3998\ : InMux
    port map (
            O => \N__17550\,
            I => \N__17544\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__17549\,
            I => \N__17541\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__17544\,
            I => \N__17538\
        );

    \I__3995\ : InMux
    port map (
            O => \N__17541\,
            I => \N__17535\
        );

    \I__3994\ : Span4Mux_v
    port map (
            O => \N__17538\,
            I => \N__17532\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__17535\,
            I => \N__17529\
        );

    \I__3992\ : Odrv4
    port map (
            O => \N__17532\,
            I => \bluejay_data_inst.n5_adj_653\
        );

    \I__3991\ : Odrv12
    port map (
            O => \N__17529\,
            I => \bluejay_data_inst.n5_adj_653\
        );

    \I__3990\ : InMux
    port map (
            O => \N__17524\,
            I => \N__17517\
        );

    \I__3989\ : InMux
    port map (
            O => \N__17523\,
            I => \N__17517\
        );

    \I__3988\ : InMux
    port map (
            O => \N__17522\,
            I => \N__17514\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__17517\,
            I => \N__17511\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__17514\,
            I => \N__17508\
        );

    \I__3985\ : Odrv12
    port map (
            O => \N__17511\,
            I => \bluejay_data_inst.n3602\
        );

    \I__3984\ : Odrv4
    port map (
            O => \N__17508\,
            I => \bluejay_data_inst.n3602\
        );

    \I__3983\ : SRMux
    port map (
            O => \N__17503\,
            I => \N__17500\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__17500\,
            I => \N__17497\
        );

    \I__3981\ : Odrv4
    port map (
            O => \N__17497\,
            I => n15
        );

    \I__3980\ : InMux
    port map (
            O => \N__17494\,
            I => \N__17489\
        );

    \I__3979\ : CascadeMux
    port map (
            O => \N__17493\,
            I => \N__17483\
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__17492\,
            I => \N__17477\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__17489\,
            I => \N__17471\
        );

    \I__3976\ : InMux
    port map (
            O => \N__17488\,
            I => \N__17468\
        );

    \I__3975\ : InMux
    port map (
            O => \N__17487\,
            I => \N__17463\
        );

    \I__3974\ : InMux
    port map (
            O => \N__17486\,
            I => \N__17463\
        );

    \I__3973\ : InMux
    port map (
            O => \N__17483\,
            I => \N__17460\
        );

    \I__3972\ : InMux
    port map (
            O => \N__17482\,
            I => \N__17457\
        );

    \I__3971\ : InMux
    port map (
            O => \N__17481\,
            I => \N__17452\
        );

    \I__3970\ : InMux
    port map (
            O => \N__17480\,
            I => \N__17452\
        );

    \I__3969\ : InMux
    port map (
            O => \N__17477\,
            I => \N__17447\
        );

    \I__3968\ : InMux
    port map (
            O => \N__17476\,
            I => \N__17447\
        );

    \I__3967\ : InMux
    port map (
            O => \N__17475\,
            I => \N__17442\
        );

    \I__3966\ : InMux
    port map (
            O => \N__17474\,
            I => \N__17442\
        );

    \I__3965\ : Span4Mux_h
    port map (
            O => \N__17471\,
            I => \N__17439\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__17468\,
            I => \N__17432\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__17463\,
            I => \N__17432\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__17460\,
            I => \N__17432\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__17457\,
            I => \bluejay_data_inst.n1394\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__17452\,
            I => \bluejay_data_inst.n1394\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__17447\,
            I => \bluejay_data_inst.n1394\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__17442\,
            I => \bluejay_data_inst.n1394\
        );

    \I__3957\ : Odrv4
    port map (
            O => \N__17439\,
            I => \bluejay_data_inst.n1394\
        );

    \I__3956\ : Odrv12
    port map (
            O => \N__17432\,
            I => \bluejay_data_inst.n1394\
        );

    \I__3955\ : InMux
    port map (
            O => \N__17419\,
            I => \N__17416\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__17416\,
            I => \N__17413\
        );

    \I__3953\ : Odrv4
    port map (
            O => \N__17413\,
            I => \bluejay_data_inst.n1133\
        );

    \I__3952\ : InMux
    port map (
            O => \N__17410\,
            I => \N__17402\
        );

    \I__3951\ : InMux
    port map (
            O => \N__17409\,
            I => \N__17402\
        );

    \I__3950\ : InMux
    port map (
            O => \N__17408\,
            I => \N__17399\
        );

    \I__3949\ : InMux
    port map (
            O => \N__17407\,
            I => \N__17395\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__17402\,
            I => \N__17392\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__17399\,
            I => \N__17389\
        );

    \I__3946\ : InMux
    port map (
            O => \N__17398\,
            I => \N__17386\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__17395\,
            I => \N__17383\
        );

    \I__3944\ : Span4Mux_h
    port map (
            O => \N__17392\,
            I => \N__17378\
        );

    \I__3943\ : Span4Mux_h
    port map (
            O => \N__17389\,
            I => \N__17378\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__17386\,
            I => \bluejay_data_inst.state_timeout_counter_5\
        );

    \I__3941\ : Odrv12
    port map (
            O => \N__17383\,
            I => \bluejay_data_inst.state_timeout_counter_5\
        );

    \I__3940\ : Odrv4
    port map (
            O => \N__17378\,
            I => \bluejay_data_inst.state_timeout_counter_5\
        );

    \I__3939\ : SRMux
    port map (
            O => \N__17371\,
            I => \N__17368\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__17368\,
            I => \N__17365\
        );

    \I__3937\ : Span4Mux_v
    port map (
            O => \N__17365\,
            I => \N__17362\
        );

    \I__3936\ : Odrv4
    port map (
            O => \N__17362\,
            I => \bluejay_data_inst.n4_adj_637\
        );

    \I__3935\ : InMux
    port map (
            O => \N__17359\,
            I => \N__17356\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__17356\,
            I => \N__17353\
        );

    \I__3933\ : Sp12to4
    port map (
            O => \N__17353\,
            I => \N__17350\
        );

    \I__3932\ : Span12Mux_v
    port map (
            O => \N__17350\,
            I => \N__17347\
        );

    \I__3931\ : Odrv12
    port map (
            O => \N__17347\,
            I => \FIFO_D4_c_4\
        );

    \I__3930\ : IoInMux
    port map (
            O => \N__17344\,
            I => \N__17341\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__17341\,
            I => \N__17338\
        );

    \I__3928\ : Span4Mux_s1_v
    port map (
            O => \N__17338\,
            I => \N__17335\
        );

    \I__3927\ : Sp12to4
    port map (
            O => \N__17335\,
            I => \N__17332\
        );

    \I__3926\ : Span12Mux_s11_h
    port map (
            O => \N__17332\,
            I => \N__17329\
        );

    \I__3925\ : Span12Mux_v
    port map (
            O => \N__17329\,
            I => \N__17326\
        );

    \I__3924\ : Odrv12
    port map (
            O => \N__17326\,
            I => \DATA4_c_4\
        );

    \I__3923\ : InMux
    port map (
            O => \N__17323\,
            I => \N__17320\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__17320\,
            I => \bluejay_data_inst.n5545\
        );

    \I__3921\ : InMux
    port map (
            O => \N__17317\,
            I => \N__17312\
        );

    \I__3920\ : InMux
    port map (
            O => \N__17316\,
            I => \N__17307\
        );

    \I__3919\ : InMux
    port map (
            O => \N__17315\,
            I => \N__17304\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__17312\,
            I => \N__17301\
        );

    \I__3917\ : InMux
    port map (
            O => \N__17311\,
            I => \N__17298\
        );

    \I__3916\ : InMux
    port map (
            O => \N__17310\,
            I => \N__17295\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__17307\,
            I => \N__17292\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__17304\,
            I => \N__17285\
        );

    \I__3913\ : Span4Mux_h
    port map (
            O => \N__17301\,
            I => \N__17285\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__17298\,
            I => \N__17285\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__17295\,
            I => \bluejay_data_inst.state_timeout_counter_1\
        );

    \I__3910\ : Odrv12
    port map (
            O => \N__17292\,
            I => \bluejay_data_inst.state_timeout_counter_1\
        );

    \I__3909\ : Odrv4
    port map (
            O => \N__17285\,
            I => \bluejay_data_inst.state_timeout_counter_1\
        );

    \I__3908\ : CascadeMux
    port map (
            O => \N__17278\,
            I => \bluejay_data_inst.n10_adj_654_cascade_\
        );

    \I__3907\ : InMux
    port map (
            O => \N__17275\,
            I => \N__17272\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__17272\,
            I => \bluejay_data_inst.n49\
        );

    \I__3905\ : CascadeMux
    port map (
            O => \N__17269\,
            I => \bluejay_data_inst.n1394_cascade_\
        );

    \I__3904\ : InMux
    port map (
            O => \N__17266\,
            I => \N__17263\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__17263\,
            I => \bluejay_data_inst.n1039\
        );

    \I__3902\ : SRMux
    port map (
            O => \N__17260\,
            I => \N__17257\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__17257\,
            I => \N__17254\
        );

    \I__3900\ : Odrv4
    port map (
            O => \N__17254\,
            I => \bluejay_data_inst.n4\
        );

    \I__3899\ : InMux
    port map (
            O => \N__17251\,
            I => \N__17240\
        );

    \I__3898\ : InMux
    port map (
            O => \N__17250\,
            I => \N__17240\
        );

    \I__3897\ : InMux
    port map (
            O => \N__17249\,
            I => \N__17240\
        );

    \I__3896\ : InMux
    port map (
            O => \N__17248\,
            I => \N__17237\
        );

    \I__3895\ : InMux
    port map (
            O => \N__17247\,
            I => \N__17234\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__17240\,
            I => \bluejay_data_inst.state_timeout_counter_4\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__17237\,
            I => \bluejay_data_inst.state_timeout_counter_4\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__17234\,
            I => \bluejay_data_inst.state_timeout_counter_4\
        );

    \I__3891\ : InMux
    port map (
            O => \N__17227\,
            I => \N__17219\
        );

    \I__3890\ : InMux
    port map (
            O => \N__17226\,
            I => \N__17219\
        );

    \I__3889\ : InMux
    port map (
            O => \N__17225\,
            I => \N__17216\
        );

    \I__3888\ : InMux
    port map (
            O => \N__17224\,
            I => \N__17213\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__17219\,
            I => \N__17209\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__17216\,
            I => \N__17204\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__17213\,
            I => \N__17204\
        );

    \I__3884\ : InMux
    port map (
            O => \N__17212\,
            I => \N__17201\
        );

    \I__3883\ : Span4Mux_v
    port map (
            O => \N__17209\,
            I => \N__17196\
        );

    \I__3882\ : Span4Mux_v
    port map (
            O => \N__17204\,
            I => \N__17196\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__17201\,
            I => \bluejay_data_inst.state_timeout_counter_3\
        );

    \I__3880\ : Odrv4
    port map (
            O => \N__17196\,
            I => \bluejay_data_inst.state_timeout_counter_3\
        );

    \I__3879\ : InMux
    port map (
            O => \N__17191\,
            I => \N__17188\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__17188\,
            I => \bluejay_data_inst.n14_adj_655\
        );

    \I__3877\ : InMux
    port map (
            O => \N__17185\,
            I => \N__17182\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__17182\,
            I => \N__17179\
        );

    \I__3875\ : Odrv4
    port map (
            O => \N__17179\,
            I => \bluejay_data_inst.n5544\
        );

    \I__3874\ : CascadeMux
    port map (
            O => \N__17176\,
            I => \bluejay_data_inst.state_timeout_counter_7_N_122_7_cascade_\
        );

    \I__3873\ : InMux
    port map (
            O => \N__17173\,
            I => \N__17170\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__17170\,
            I => \bluejay_data_inst.state_timeout_counter_7_N_122_7\
        );

    \I__3871\ : CascadeMux
    port map (
            O => \N__17167\,
            I => \bluejay_data_inst.n8_adj_640_cascade_\
        );

    \I__3870\ : InMux
    port map (
            O => \N__17164\,
            I => \N__17161\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__17161\,
            I => \N__17158\
        );

    \I__3868\ : Span4Mux_h
    port map (
            O => \N__17158\,
            I => \N__17155\
        );

    \I__3867\ : Odrv4
    port map (
            O => \N__17155\,
            I => \bluejay_data_inst.n51\
        );

    \I__3866\ : InMux
    port map (
            O => \N__17152\,
            I => \bluejay_data_inst.n4817\
        );

    \I__3865\ : InMux
    port map (
            O => \N__17149\,
            I => \N__17146\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__17146\,
            I => \N__17143\
        );

    \I__3863\ : Span4Mux_h
    port map (
            O => \N__17143\,
            I => \N__17140\
        );

    \I__3862\ : Odrv4
    port map (
            O => \N__17140\,
            I => \bluejay_data_inst.n50\
        );

    \I__3861\ : InMux
    port map (
            O => \N__17137\,
            I => \bluejay_data_inst.n4818\
        );

    \I__3860\ : InMux
    port map (
            O => \N__17134\,
            I => \bluejay_data_inst.n4819\
        );

    \I__3859\ : InMux
    port map (
            O => \N__17131\,
            I => \N__17128\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__17128\,
            I => \bluejay_data_inst.n48\
        );

    \I__3857\ : InMux
    port map (
            O => \N__17125\,
            I => \bluejay_data_inst.n4820\
        );

    \I__3856\ : InMux
    port map (
            O => \N__17122\,
            I => \bluejay_data_inst.n4821\
        );

    \I__3855\ : IoInMux
    port map (
            O => \N__17119\,
            I => \N__17116\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__17116\,
            I => \N__17109\
        );

    \I__3853\ : IoInMux
    port map (
            O => \N__17115\,
            I => \N__17106\
        );

    \I__3852\ : CascadeMux
    port map (
            O => \N__17114\,
            I => \N__17101\
        );

    \I__3851\ : CascadeMux
    port map (
            O => \N__17113\,
            I => \N__17097\
        );

    \I__3850\ : CascadeMux
    port map (
            O => \N__17112\,
            I => \N__17093\
        );

    \I__3849\ : IoSpan4Mux
    port map (
            O => \N__17109\,
            I => \N__17090\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__17106\,
            I => \N__17087\
        );

    \I__3847\ : InMux
    port map (
            O => \N__17105\,
            I => \N__17072\
        );

    \I__3846\ : InMux
    port map (
            O => \N__17104\,
            I => \N__17072\
        );

    \I__3845\ : InMux
    port map (
            O => \N__17101\,
            I => \N__17072\
        );

    \I__3844\ : InMux
    port map (
            O => \N__17100\,
            I => \N__17072\
        );

    \I__3843\ : InMux
    port map (
            O => \N__17097\,
            I => \N__17072\
        );

    \I__3842\ : InMux
    port map (
            O => \N__17096\,
            I => \N__17072\
        );

    \I__3841\ : InMux
    port map (
            O => \N__17093\,
            I => \N__17072\
        );

    \I__3840\ : Span4Mux_s3_h
    port map (
            O => \N__17090\,
            I => \N__17067\
        );

    \I__3839\ : Span4Mux_s3_h
    port map (
            O => \N__17087\,
            I => \N__17067\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__17072\,
            I => \N__17064\
        );

    \I__3837\ : Span4Mux_v
    port map (
            O => \N__17067\,
            I => \N__17058\
        );

    \I__3836\ : Span4Mux_v
    port map (
            O => \N__17064\,
            I => \N__17052\
        );

    \I__3835\ : CascadeMux
    port map (
            O => \N__17063\,
            I => \N__17049\
        );

    \I__3834\ : CascadeMux
    port map (
            O => \N__17062\,
            I => \N__17046\
        );

    \I__3833\ : CascadeMux
    port map (
            O => \N__17061\,
            I => \N__17043\
        );

    \I__3832\ : Sp12to4
    port map (
            O => \N__17058\,
            I => \N__17031\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__17057\,
            I => \N__17027\
        );

    \I__3830\ : CascadeMux
    port map (
            O => \N__17056\,
            I => \N__17024\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__17055\,
            I => \N__17021\
        );

    \I__3828\ : Span4Mux_h
    port map (
            O => \N__17052\,
            I => \N__17018\
        );

    \I__3827\ : InMux
    port map (
            O => \N__17049\,
            I => \N__17011\
        );

    \I__3826\ : InMux
    port map (
            O => \N__17046\,
            I => \N__17011\
        );

    \I__3825\ : InMux
    port map (
            O => \N__17043\,
            I => \N__17011\
        );

    \I__3824\ : CascadeMux
    port map (
            O => \N__17042\,
            I => \N__17008\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__17041\,
            I => \N__17005\
        );

    \I__3822\ : CascadeMux
    port map (
            O => \N__17040\,
            I => \N__16998\
        );

    \I__3821\ : CascadeMux
    port map (
            O => \N__17039\,
            I => \N__16994\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__17038\,
            I => \N__16991\
        );

    \I__3819\ : CascadeMux
    port map (
            O => \N__17037\,
            I => \N__16988\
        );

    \I__3818\ : CascadeMux
    port map (
            O => \N__17036\,
            I => \N__16985\
        );

    \I__3817\ : CascadeMux
    port map (
            O => \N__17035\,
            I => \N__16982\
        );

    \I__3816\ : CascadeMux
    port map (
            O => \N__17034\,
            I => \N__16979\
        );

    \I__3815\ : Span12Mux_h
    port map (
            O => \N__17031\,
            I => \N__16976\
        );

    \I__3814\ : InMux
    port map (
            O => \N__17030\,
            I => \N__16967\
        );

    \I__3813\ : InMux
    port map (
            O => \N__17027\,
            I => \N__16967\
        );

    \I__3812\ : InMux
    port map (
            O => \N__17024\,
            I => \N__16967\
        );

    \I__3811\ : InMux
    port map (
            O => \N__17021\,
            I => \N__16967\
        );

    \I__3810\ : Span4Mux_h
    port map (
            O => \N__17018\,
            I => \N__16962\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__17011\,
            I => \N__16962\
        );

    \I__3808\ : InMux
    port map (
            O => \N__17008\,
            I => \N__16947\
        );

    \I__3807\ : InMux
    port map (
            O => \N__17005\,
            I => \N__16947\
        );

    \I__3806\ : InMux
    port map (
            O => \N__17004\,
            I => \N__16947\
        );

    \I__3805\ : InMux
    port map (
            O => \N__17003\,
            I => \N__16947\
        );

    \I__3804\ : InMux
    port map (
            O => \N__17002\,
            I => \N__16947\
        );

    \I__3803\ : InMux
    port map (
            O => \N__17001\,
            I => \N__16947\
        );

    \I__3802\ : InMux
    port map (
            O => \N__16998\,
            I => \N__16947\
        );

    \I__3801\ : InMux
    port map (
            O => \N__16997\,
            I => \N__16938\
        );

    \I__3800\ : InMux
    port map (
            O => \N__16994\,
            I => \N__16938\
        );

    \I__3799\ : InMux
    port map (
            O => \N__16991\,
            I => \N__16938\
        );

    \I__3798\ : InMux
    port map (
            O => \N__16988\,
            I => \N__16938\
        );

    \I__3797\ : InMux
    port map (
            O => \N__16985\,
            I => \N__16931\
        );

    \I__3796\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16931\
        );

    \I__3795\ : InMux
    port map (
            O => \N__16979\,
            I => \N__16931\
        );

    \I__3794\ : Span12Mux_v
    port map (
            O => \N__16976\,
            I => \N__16928\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__16967\,
            I => \N__16925\
        );

    \I__3792\ : Span4Mux_v
    port map (
            O => \N__16962\,
            I => \N__16920\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__16947\,
            I => \N__16920\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__16938\,
            I => \N__16915\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__16931\,
            I => \N__16915\
        );

    \I__3788\ : Odrv12
    port map (
            O => \N__16928\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3787\ : Odrv12
    port map (
            O => \N__16925\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__16920\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3785\ : Odrv4
    port map (
            O => \N__16915\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3784\ : InMux
    port map (
            O => \N__16906\,
            I => \bluejay_data_inst.n4822\
        );

    \I__3783\ : CascadeMux
    port map (
            O => \N__16903\,
            I => \bluejay_data_inst.state_timeout_counter_7_N_122_4_cascade_\
        );

    \I__3782\ : InMux
    port map (
            O => \N__16900\,
            I => \N__16897\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__16897\,
            I => \bluejay_data_inst.state_timeout_counter_7_N_122_4\
        );

    \I__3780\ : CascadeMux
    port map (
            O => \N__16894\,
            I => \bluejay_data_inst.n8_cascade_\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__16891\,
            I => \N__16888\
        );

    \I__3778\ : InMux
    port map (
            O => \N__16888\,
            I => \N__16885\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__16885\,
            I => \N__16881\
        );

    \I__3776\ : InMux
    port map (
            O => \N__16884\,
            I => \N__16878\
        );

    \I__3775\ : Odrv4
    port map (
            O => \N__16881\,
            I => \bluejay_data_inst.h_counter_2\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__16878\,
            I => \bluejay_data_inst.h_counter_2\
        );

    \I__3773\ : InMux
    port map (
            O => \N__16873\,
            I => \bluejay_data_inst.n4859\
        );

    \I__3772\ : InMux
    port map (
            O => \N__16870\,
            I => \N__16866\
        );

    \I__3771\ : InMux
    port map (
            O => \N__16869\,
            I => \N__16863\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__16866\,
            I => \bluejay_data_inst.h_counter_3\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__16863\,
            I => \bluejay_data_inst.h_counter_3\
        );

    \I__3768\ : InMux
    port map (
            O => \N__16858\,
            I => \N__16855\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__16855\,
            I => \bluejay_data_inst.n5547\
        );

    \I__3766\ : InMux
    port map (
            O => \N__16852\,
            I => \bluejay_data_inst.n4860\
        );

    \I__3765\ : CascadeMux
    port map (
            O => \N__16849\,
            I => \N__16846\
        );

    \I__3764\ : InMux
    port map (
            O => \N__16846\,
            I => \N__16842\
        );

    \I__3763\ : InMux
    port map (
            O => \N__16845\,
            I => \N__16839\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__16842\,
            I => \bluejay_data_inst.h_counter_4\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__16839\,
            I => \bluejay_data_inst.h_counter_4\
        );

    \I__3760\ : InMux
    port map (
            O => \N__16834\,
            I => \bluejay_data_inst.n4861\
        );

    \I__3759\ : InMux
    port map (
            O => \N__16831\,
            I => \N__16823\
        );

    \I__3758\ : InMux
    port map (
            O => \N__16830\,
            I => \N__16823\
        );

    \I__3757\ : InMux
    port map (
            O => \N__16829\,
            I => \N__16818\
        );

    \I__3756\ : InMux
    port map (
            O => \N__16828\,
            I => \N__16812\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__16823\,
            I => \N__16809\
        );

    \I__3754\ : InMux
    port map (
            O => \N__16822\,
            I => \N__16804\
        );

    \I__3753\ : InMux
    port map (
            O => \N__16821\,
            I => \N__16804\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__16818\,
            I => \N__16801\
        );

    \I__3751\ : InMux
    port map (
            O => \N__16817\,
            I => \N__16796\
        );

    \I__3750\ : InMux
    port map (
            O => \N__16816\,
            I => \N__16796\
        );

    \I__3749\ : InMux
    port map (
            O => \N__16815\,
            I => \N__16793\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__16812\,
            I => \N__16790\
        );

    \I__3747\ : Odrv12
    port map (
            O => \N__16809\,
            I => \bluejay_data_inst.valid_o_N_155\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__16804\,
            I => \bluejay_data_inst.valid_o_N_155\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__16801\,
            I => \bluejay_data_inst.valid_o_N_155\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__16796\,
            I => \bluejay_data_inst.valid_o_N_155\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__16793\,
            I => \bluejay_data_inst.valid_o_N_155\
        );

    \I__3742\ : Odrv4
    port map (
            O => \N__16790\,
            I => \bluejay_data_inst.valid_o_N_155\
        );

    \I__3741\ : InMux
    port map (
            O => \N__16777\,
            I => \N__16773\
        );

    \I__3740\ : InMux
    port map (
            O => \N__16776\,
            I => \N__16770\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__16773\,
            I => \bluejay_data_inst.h_counter_5\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__16770\,
            I => \bluejay_data_inst.h_counter_5\
        );

    \I__3737\ : InMux
    port map (
            O => \N__16765\,
            I => \N__16762\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__16762\,
            I => \bluejay_data_inst.n5548\
        );

    \I__3735\ : InMux
    port map (
            O => \N__16759\,
            I => \bluejay_data_inst.n4862\
        );

    \I__3734\ : CascadeMux
    port map (
            O => \N__16756\,
            I => \N__16753\
        );

    \I__3733\ : InMux
    port map (
            O => \N__16753\,
            I => \N__16749\
        );

    \I__3732\ : InMux
    port map (
            O => \N__16752\,
            I => \N__16746\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__16749\,
            I => \bluejay_data_inst.h_counter_6\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__16746\,
            I => \bluejay_data_inst.h_counter_6\
        );

    \I__3729\ : InMux
    port map (
            O => \N__16741\,
            I => \bluejay_data_inst.n4863\
        );

    \I__3728\ : InMux
    port map (
            O => \N__16738\,
            I => \bluejay_data_inst.n4864\
        );

    \I__3727\ : CascadeMux
    port map (
            O => \N__16735\,
            I => \N__16732\
        );

    \I__3726\ : InMux
    port map (
            O => \N__16732\,
            I => \N__16728\
        );

    \I__3725\ : InMux
    port map (
            O => \N__16731\,
            I => \N__16725\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__16728\,
            I => \N__16722\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__16725\,
            I => \bluejay_data_inst.h_counter_7\
        );

    \I__3722\ : Odrv4
    port map (
            O => \N__16722\,
            I => \bluejay_data_inst.h_counter_7\
        );

    \I__3721\ : CEMux
    port map (
            O => \N__16717\,
            I => \N__16713\
        );

    \I__3720\ : CEMux
    port map (
            O => \N__16716\,
            I => \N__16710\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__16713\,
            I => \N__16707\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__16710\,
            I => \N__16704\
        );

    \I__3717\ : Span4Mux_h
    port map (
            O => \N__16707\,
            I => \N__16699\
        );

    \I__3716\ : Span4Mux_h
    port map (
            O => \N__16704\,
            I => \N__16699\
        );

    \I__3715\ : Span4Mux_h
    port map (
            O => \N__16699\,
            I => \N__16695\
        );

    \I__3714\ : InMux
    port map (
            O => \N__16698\,
            I => \N__16692\
        );

    \I__3713\ : Odrv4
    port map (
            O => \N__16695\,
            I => n2555
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__16692\,
            I => n2555
        );

    \I__3711\ : SRMux
    port map (
            O => \N__16687\,
            I => \N__16684\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__16684\,
            I => \N__16681\
        );

    \I__3709\ : Span4Mux_h
    port map (
            O => \N__16681\,
            I => \N__16678\
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__16678\,
            I => \bluejay_data_inst.n2693\
        );

    \I__3707\ : InMux
    port map (
            O => \N__16675\,
            I => \bfn_17_8_0_\
        );

    \I__3706\ : InMux
    port map (
            O => \N__16672\,
            I => \N__16669\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__16669\,
            I => \bluejay_data_inst.n5527\
        );

    \I__3704\ : InMux
    port map (
            O => \N__16666\,
            I => \bluejay_data_inst.n4816\
        );

    \I__3703\ : CascadeMux
    port map (
            O => \N__16663\,
            I => \N__16653\
        );

    \I__3702\ : CascadeMux
    port map (
            O => \N__16662\,
            I => \N__16646\
        );

    \I__3701\ : InMux
    port map (
            O => \N__16661\,
            I => \N__16635\
        );

    \I__3700\ : InMux
    port map (
            O => \N__16660\,
            I => \N__16635\
        );

    \I__3699\ : InMux
    port map (
            O => \N__16659\,
            I => \N__16618\
        );

    \I__3698\ : InMux
    port map (
            O => \N__16658\,
            I => \N__16618\
        );

    \I__3697\ : InMux
    port map (
            O => \N__16657\,
            I => \N__16618\
        );

    \I__3696\ : InMux
    port map (
            O => \N__16656\,
            I => \N__16618\
        );

    \I__3695\ : InMux
    port map (
            O => \N__16653\,
            I => \N__16618\
        );

    \I__3694\ : InMux
    port map (
            O => \N__16652\,
            I => \N__16618\
        );

    \I__3693\ : InMux
    port map (
            O => \N__16651\,
            I => \N__16618\
        );

    \I__3692\ : InMux
    port map (
            O => \N__16650\,
            I => \N__16618\
        );

    \I__3691\ : InMux
    port map (
            O => \N__16649\,
            I => \N__16611\
        );

    \I__3690\ : InMux
    port map (
            O => \N__16646\,
            I => \N__16611\
        );

    \I__3689\ : InMux
    port map (
            O => \N__16645\,
            I => \N__16611\
        );

    \I__3688\ : InMux
    port map (
            O => \N__16644\,
            I => \N__16606\
        );

    \I__3687\ : InMux
    port map (
            O => \N__16643\,
            I => \N__16606\
        );

    \I__3686\ : InMux
    port map (
            O => \N__16642\,
            I => \N__16603\
        );

    \I__3685\ : InMux
    port map (
            O => \N__16641\,
            I => \N__16600\
        );

    \I__3684\ : InMux
    port map (
            O => \N__16640\,
            I => \N__16597\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__16635\,
            I => n5
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__16618\,
            I => n5
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__16611\,
            I => n5
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__16606\,
            I => n5
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__16603\,
            I => n5
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__16600\,
            I => n5
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__16597\,
            I => n5
        );

    \I__3676\ : CascadeMux
    port map (
            O => \N__16582\,
            I => \bluejay_data_inst.n3631_cascade_\
        );

    \I__3675\ : SRMux
    port map (
            O => \N__16579\,
            I => \N__16569\
        );

    \I__3674\ : SRMux
    port map (
            O => \N__16578\,
            I => \N__16562\
        );

    \I__3673\ : SRMux
    port map (
            O => \N__16577\,
            I => \N__16559\
        );

    \I__3672\ : InMux
    port map (
            O => \N__16576\,
            I => \N__16554\
        );

    \I__3671\ : InMux
    port map (
            O => \N__16575\,
            I => \N__16551\
        );

    \I__3670\ : InMux
    port map (
            O => \N__16574\,
            I => \N__16548\
        );

    \I__3669\ : SRMux
    port map (
            O => \N__16573\,
            I => \N__16540\
        );

    \I__3668\ : InMux
    port map (
            O => \N__16572\,
            I => \N__16537\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__16569\,
            I => \N__16534\
        );

    \I__3666\ : SRMux
    port map (
            O => \N__16568\,
            I => \N__16531\
        );

    \I__3665\ : SRMux
    port map (
            O => \N__16567\,
            I => \N__16528\
        );

    \I__3664\ : InMux
    port map (
            O => \N__16566\,
            I => \N__16525\
        );

    \I__3663\ : SRMux
    port map (
            O => \N__16565\,
            I => \N__16520\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__16562\,
            I => \N__16517\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__16559\,
            I => \N__16514\
        );

    \I__3660\ : SRMux
    port map (
            O => \N__16558\,
            I => \N__16511\
        );

    \I__3659\ : CascadeMux
    port map (
            O => \N__16557\,
            I => \N__16508\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__16554\,
            I => \N__16504\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__16551\,
            I => \N__16499\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__16548\,
            I => \N__16499\
        );

    \I__3655\ : InMux
    port map (
            O => \N__16547\,
            I => \N__16494\
        );

    \I__3654\ : InMux
    port map (
            O => \N__16546\,
            I => \N__16494\
        );

    \I__3653\ : SRMux
    port map (
            O => \N__16545\,
            I => \N__16489\
        );

    \I__3652\ : SRMux
    port map (
            O => \N__16544\,
            I => \N__16486\
        );

    \I__3651\ : SRMux
    port map (
            O => \N__16543\,
            I => \N__16483\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__16540\,
            I => \N__16480\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__16537\,
            I => \N__16476\
        );

    \I__3648\ : Span4Mux_h
    port map (
            O => \N__16534\,
            I => \N__16467\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__16531\,
            I => \N__16467\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__16528\,
            I => \N__16467\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__16525\,
            I => \N__16467\
        );

    \I__3644\ : InMux
    port map (
            O => \N__16524\,
            I => \N__16464\
        );

    \I__3643\ : SRMux
    port map (
            O => \N__16523\,
            I => \N__16461\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__16520\,
            I => \N__16458\
        );

    \I__3641\ : Span4Mux_v
    port map (
            O => \N__16517\,
            I => \N__16451\
        );

    \I__3640\ : Span4Mux_h
    port map (
            O => \N__16514\,
            I => \N__16451\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__16511\,
            I => \N__16451\
        );

    \I__3638\ : InMux
    port map (
            O => \N__16508\,
            I => \N__16446\
        );

    \I__3637\ : InMux
    port map (
            O => \N__16507\,
            I => \N__16446\
        );

    \I__3636\ : Span4Mux_h
    port map (
            O => \N__16504\,
            I => \N__16439\
        );

    \I__3635\ : Span4Mux_v
    port map (
            O => \N__16499\,
            I => \N__16439\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__16494\,
            I => \N__16439\
        );

    \I__3633\ : InMux
    port map (
            O => \N__16493\,
            I => \N__16436\
        );

    \I__3632\ : InMux
    port map (
            O => \N__16492\,
            I => \N__16431\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__16489\,
            I => \N__16428\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__16486\,
            I => \N__16422\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__16483\,
            I => \N__16422\
        );

    \I__3628\ : Span4Mux_v
    port map (
            O => \N__16480\,
            I => \N__16419\
        );

    \I__3627\ : InMux
    port map (
            O => \N__16479\,
            I => \N__16416\
        );

    \I__3626\ : Span4Mux_v
    port map (
            O => \N__16476\,
            I => \N__16407\
        );

    \I__3625\ : Span4Mux_v
    port map (
            O => \N__16467\,
            I => \N__16407\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__16464\,
            I => \N__16404\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__16461\,
            I => \N__16400\
        );

    \I__3622\ : Span4Mux_v
    port map (
            O => \N__16458\,
            I => \N__16395\
        );

    \I__3621\ : Span4Mux_h
    port map (
            O => \N__16451\,
            I => \N__16395\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__16446\,
            I => \N__16388\
        );

    \I__3619\ : Span4Mux_h
    port map (
            O => \N__16439\,
            I => \N__16388\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__16436\,
            I => \N__16388\
        );

    \I__3617\ : InMux
    port map (
            O => \N__16435\,
            I => \N__16383\
        );

    \I__3616\ : InMux
    port map (
            O => \N__16434\,
            I => \N__16383\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__16431\,
            I => \N__16380\
        );

    \I__3614\ : Span4Mux_v
    port map (
            O => \N__16428\,
            I => \N__16377\
        );

    \I__3613\ : InMux
    port map (
            O => \N__16427\,
            I => \N__16374\
        );

    \I__3612\ : Span4Mux_h
    port map (
            O => \N__16422\,
            I => \N__16367\
        );

    \I__3611\ : Span4Mux_h
    port map (
            O => \N__16419\,
            I => \N__16367\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__16416\,
            I => \N__16367\
        );

    \I__3609\ : InMux
    port map (
            O => \N__16415\,
            I => \N__16364\
        );

    \I__3608\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16361\
        );

    \I__3607\ : InMux
    port map (
            O => \N__16413\,
            I => \N__16356\
        );

    \I__3606\ : InMux
    port map (
            O => \N__16412\,
            I => \N__16356\
        );

    \I__3605\ : Sp12to4
    port map (
            O => \N__16407\,
            I => \N__16351\
        );

    \I__3604\ : Span12Mux_v
    port map (
            O => \N__16404\,
            I => \N__16351\
        );

    \I__3603\ : InMux
    port map (
            O => \N__16403\,
            I => \N__16348\
        );

    \I__3602\ : Span4Mux_v
    port map (
            O => \N__16400\,
            I => \N__16337\
        );

    \I__3601\ : Span4Mux_h
    port map (
            O => \N__16395\,
            I => \N__16337\
        );

    \I__3600\ : Span4Mux_v
    port map (
            O => \N__16388\,
            I => \N__16337\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__16383\,
            I => \N__16337\
        );

    \I__3598\ : Span4Mux_h
    port map (
            O => \N__16380\,
            I => \N__16337\
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__16377\,
            I => reset_all_w
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__16374\,
            I => reset_all_w
        );

    \I__3595\ : Odrv4
    port map (
            O => \N__16367\,
            I => reset_all_w
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__16364\,
            I => reset_all_w
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__16361\,
            I => reset_all_w
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__16356\,
            I => reset_all_w
        );

    \I__3591\ : Odrv12
    port map (
            O => \N__16351\,
            I => reset_all_w
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__16348\,
            I => reset_all_w
        );

    \I__3589\ : Odrv4
    port map (
            O => \N__16337\,
            I => reset_all_w
        );

    \I__3588\ : InMux
    port map (
            O => \N__16318\,
            I => \N__16315\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__16315\,
            I => \N__16312\
        );

    \I__3586\ : Odrv12
    port map (
            O => \N__16312\,
            I => \bluejay_data_inst.state_timeout_counter_7_N_122_5\
        );

    \I__3585\ : InMux
    port map (
            O => \N__16309\,
            I => \N__16306\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__16306\,
            I => \N__16303\
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__16303\,
            I => \bluejay_data_inst.n4266\
        );

    \I__3582\ : SRMux
    port map (
            O => \N__16300\,
            I => \N__16297\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__16297\,
            I => \N__16294\
        );

    \I__3580\ : Odrv12
    port map (
            O => \N__16294\,
            I => \bluejay_data_inst.n4_adj_652\
        );

    \I__3579\ : InMux
    port map (
            O => \N__16291\,
            I => \N__16288\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__16288\,
            I => \N__16285\
        );

    \I__3577\ : Span4Mux_v
    port map (
            O => \N__16285\,
            I => \N__16282\
        );

    \I__3576\ : Sp12to4
    port map (
            O => \N__16282\,
            I => \N__16279\
        );

    \I__3575\ : Span12Mux_h
    port map (
            O => \N__16279\,
            I => \N__16276\
        );

    \I__3574\ : Span12Mux_v
    port map (
            O => \N__16276\,
            I => \N__16273\
        );

    \I__3573\ : Odrv12
    port map (
            O => \N__16273\,
            I => \FIFO_D0_c_0\
        );

    \I__3572\ : IoInMux
    port map (
            O => \N__16270\,
            I => \N__16267\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__16267\,
            I => \N__16264\
        );

    \I__3570\ : IoSpan4Mux
    port map (
            O => \N__16264\,
            I => \N__16261\
        );

    \I__3569\ : Sp12to4
    port map (
            O => \N__16261\,
            I => \N__16258\
        );

    \I__3568\ : Span12Mux_v
    port map (
            O => \N__16258\,
            I => \N__16255\
        );

    \I__3567\ : Span12Mux_h
    port map (
            O => \N__16255\,
            I => \N__16252\
        );

    \I__3566\ : Odrv12
    port map (
            O => \N__16252\,
            I => \DATA0_c_0\
        );

    \I__3565\ : IoInMux
    port map (
            O => \N__16249\,
            I => \N__16246\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__16246\,
            I => \N__16243\
        );

    \I__3563\ : IoSpan4Mux
    port map (
            O => \N__16243\,
            I => \N__16240\
        );

    \I__3562\ : Span4Mux_s3_h
    port map (
            O => \N__16240\,
            I => \N__16236\
        );

    \I__3561\ : InMux
    port map (
            O => \N__16239\,
            I => \N__16233\
        );

    \I__3560\ : Span4Mux_v
    port map (
            O => \N__16236\,
            I => \N__16230\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__16233\,
            I => \N__16227\
        );

    \I__3558\ : Sp12to4
    port map (
            O => \N__16230\,
            I => \N__16224\
        );

    \I__3557\ : Span4Mux_v
    port map (
            O => \N__16227\,
            I => \N__16221\
        );

    \I__3556\ : Span12Mux_h
    port map (
            O => \N__16224\,
            I => \N__16216\
        );

    \I__3555\ : Sp12to4
    port map (
            O => \N__16221\,
            I => \N__16216\
        );

    \I__3554\ : Span12Mux_h
    port map (
            O => \N__16216\,
            I => \N__16213\
        );

    \I__3553\ : Odrv12
    port map (
            O => \N__16213\,
            I => \DEBUG_6_c_22_c\
        );

    \I__3552\ : IoInMux
    port map (
            O => \N__16210\,
            I => \N__16207\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__16207\,
            I => \N__16204\
        );

    \I__3550\ : Span4Mux_s3_v
    port map (
            O => \N__16204\,
            I => \N__16201\
        );

    \I__3549\ : Sp12to4
    port map (
            O => \N__16201\,
            I => \N__16197\
        );

    \I__3548\ : IoInMux
    port map (
            O => \N__16200\,
            I => \N__16194\
        );

    \I__3547\ : Span12Mux_s11_h
    port map (
            O => \N__16197\,
            I => \N__16191\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__16194\,
            I => \N__16188\
        );

    \I__3545\ : Span12Mux_v
    port map (
            O => \N__16191\,
            I => \N__16183\
        );

    \I__3544\ : Span12Mux_s11_h
    port map (
            O => \N__16188\,
            I => \N__16183\
        );

    \I__3543\ : Odrv12
    port map (
            O => \N__16183\,
            I => \DEBUG_5_c\
        );

    \I__3542\ : SRMux
    port map (
            O => \N__16180\,
            I => \N__16174\
        );

    \I__3541\ : SRMux
    port map (
            O => \N__16179\,
            I => \N__16171\
        );

    \I__3540\ : InMux
    port map (
            O => \N__16178\,
            I => \N__16168\
        );

    \I__3539\ : InMux
    port map (
            O => \N__16177\,
            I => \N__16165\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__16174\,
            I => \N__16162\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__16171\,
            I => \N__16159\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__16168\,
            I => \N__16156\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__16165\,
            I => \N__16153\
        );

    \I__3534\ : Span4Mux_h
    port map (
            O => \N__16162\,
            I => \N__16148\
        );

    \I__3533\ : Span4Mux_h
    port map (
            O => \N__16159\,
            I => \N__16144\
        );

    \I__3532\ : Span4Mux_h
    port map (
            O => \N__16156\,
            I => \N__16141\
        );

    \I__3531\ : Span4Mux_h
    port map (
            O => \N__16153\,
            I => \N__16137\
        );

    \I__3530\ : InMux
    port map (
            O => \N__16152\,
            I => \N__16134\
        );

    \I__3529\ : InMux
    port map (
            O => \N__16151\,
            I => \N__16131\
        );

    \I__3528\ : Sp12to4
    port map (
            O => \N__16148\,
            I => \N__16128\
        );

    \I__3527\ : InMux
    port map (
            O => \N__16147\,
            I => \N__16125\
        );

    \I__3526\ : Span4Mux_h
    port map (
            O => \N__16144\,
            I => \N__16120\
        );

    \I__3525\ : Span4Mux_h
    port map (
            O => \N__16141\,
            I => \N__16120\
        );

    \I__3524\ : InMux
    port map (
            O => \N__16140\,
            I => \N__16117\
        );

    \I__3523\ : Span4Mux_h
    port map (
            O => \N__16137\,
            I => \N__16114\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__16134\,
            I => \N__16109\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__16131\,
            I => \N__16109\
        );

    \I__3520\ : Odrv12
    port map (
            O => \N__16128\,
            I => \r_SM_Main_2_adj_659\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__16125\,
            I => \r_SM_Main_2_adj_659\
        );

    \I__3518\ : Odrv4
    port map (
            O => \N__16120\,
            I => \r_SM_Main_2_adj_659\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__16117\,
            I => \r_SM_Main_2_adj_659\
        );

    \I__3516\ : Odrv4
    port map (
            O => \N__16114\,
            I => \r_SM_Main_2_adj_659\
        );

    \I__3515\ : Odrv12
    port map (
            O => \N__16109\,
            I => \r_SM_Main_2_adj_659\
        );

    \I__3514\ : CEMux
    port map (
            O => \N__16096\,
            I => \N__16091\
        );

    \I__3513\ : CEMux
    port map (
            O => \N__16095\,
            I => \N__16088\
        );

    \I__3512\ : CEMux
    port map (
            O => \N__16094\,
            I => \N__16085\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__16091\,
            I => \N__16082\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__16088\,
            I => \N__16079\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__16085\,
            I => \N__16076\
        );

    \I__3508\ : Span4Mux_s1_h
    port map (
            O => \N__16082\,
            I => \N__16073\
        );

    \I__3507\ : Span4Mux_h
    port map (
            O => \N__16079\,
            I => \N__16070\
        );

    \I__3506\ : Sp12to4
    port map (
            O => \N__16076\,
            I => \N__16067\
        );

    \I__3505\ : Sp12to4
    port map (
            O => \N__16073\,
            I => \N__16064\
        );

    \I__3504\ : Span4Mux_h
    port map (
            O => \N__16070\,
            I => \N__16061\
        );

    \I__3503\ : Span12Mux_h
    port map (
            O => \N__16067\,
            I => \N__16056\
        );

    \I__3502\ : Span12Mux_s11_v
    port map (
            O => \N__16064\,
            I => \N__16056\
        );

    \I__3501\ : Odrv4
    port map (
            O => \N__16061\,
            I => \pc_tx.n1\
        );

    \I__3500\ : Odrv12
    port map (
            O => \N__16056\,
            I => \pc_tx.n1\
        );

    \I__3499\ : InMux
    port map (
            O => \N__16051\,
            I => \N__16047\
        );

    \I__3498\ : InMux
    port map (
            O => \N__16050\,
            I => \N__16044\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__16047\,
            I => \N__16041\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__16044\,
            I => \bluejay_data_inst.h_counter_0\
        );

    \I__3495\ : Odrv4
    port map (
            O => \N__16041\,
            I => \bluejay_data_inst.h_counter_0\
        );

    \I__3494\ : InMux
    port map (
            O => \N__16036\,
            I => \bfn_17_7_0_\
        );

    \I__3493\ : InMux
    port map (
            O => \N__16033\,
            I => \N__16029\
        );

    \I__3492\ : InMux
    port map (
            O => \N__16032\,
            I => \N__16026\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__16029\,
            I => \N__16023\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__16026\,
            I => \N__16018\
        );

    \I__3489\ : Span4Mux_h
    port map (
            O => \N__16023\,
            I => \N__16018\
        );

    \I__3488\ : Odrv4
    port map (
            O => \N__16018\,
            I => \bluejay_data_inst.h_counter_1\
        );

    \I__3487\ : InMux
    port map (
            O => \N__16015\,
            I => \bluejay_data_inst.n4858\
        );

    \I__3486\ : InMux
    port map (
            O => \N__16012\,
            I => \N__16009\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__16009\,
            I => \bluejay_data_inst.n31\
        );

    \I__3484\ : CascadeMux
    port map (
            O => \N__16006\,
            I => \bluejay_data_inst.state_timeout_counter_7_N_122_5_cascade_\
        );

    \I__3483\ : IoInMux
    port map (
            O => \N__16003\,
            I => \N__16000\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__16000\,
            I => \N__15997\
        );

    \I__3481\ : Span4Mux_s3_h
    port map (
            O => \N__15997\,
            I => \N__15993\
        );

    \I__3480\ : CascadeMux
    port map (
            O => \N__15996\,
            I => \N__15990\
        );

    \I__3479\ : Span4Mux_h
    port map (
            O => \N__15993\,
            I => \N__15987\
        );

    \I__3478\ : InMux
    port map (
            O => \N__15990\,
            I => \N__15984\
        );

    \I__3477\ : Span4Mux_h
    port map (
            O => \N__15987\,
            I => \N__15980\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__15984\,
            I => \N__15977\
        );

    \I__3475\ : InMux
    port map (
            O => \N__15983\,
            I => \N__15974\
        );

    \I__3474\ : Odrv4
    port map (
            O => \N__15980\,
            I => \DEBUG_3_c\
        );

    \I__3473\ : Odrv12
    port map (
            O => \N__15977\,
            I => \DEBUG_3_c\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__15974\,
            I => \DEBUG_3_c\
        );

    \I__3471\ : InMux
    port map (
            O => \N__15967\,
            I => \N__15964\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__15964\,
            I => \bluejay_data_inst.n11\
        );

    \I__3469\ : InMux
    port map (
            O => \N__15961\,
            I => \N__15958\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__15958\,
            I => \bluejay_data_inst.n9\
        );

    \I__3467\ : InMux
    port map (
            O => \N__15955\,
            I => \N__15949\
        );

    \I__3466\ : InMux
    port map (
            O => \N__15954\,
            I => \N__15949\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__15949\,
            I => \bluejay_data_inst.n4252\
        );

    \I__3464\ : SRMux
    port map (
            O => \N__15946\,
            I => \N__15943\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__15943\,
            I => \N__15940\
        );

    \I__3462\ : Span4Mux_v
    port map (
            O => \N__15940\,
            I => \N__15937\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__15937\,
            I => \bluejay_data_inst.n4_adj_648\
        );

    \I__3460\ : CascadeMux
    port map (
            O => \N__15934\,
            I => \bluejay_data_inst.n3627_cascade_\
        );

    \I__3459\ : IoInMux
    port map (
            O => \N__15931\,
            I => \N__15928\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__15928\,
            I => \N__15924\
        );

    \I__3457\ : CascadeMux
    port map (
            O => \N__15927\,
            I => \N__15920\
        );

    \I__3456\ : Span12Mux_s5_h
    port map (
            O => \N__15924\,
            I => \N__15917\
        );

    \I__3455\ : InMux
    port map (
            O => \N__15923\,
            I => \N__15914\
        );

    \I__3454\ : InMux
    port map (
            O => \N__15920\,
            I => \N__15911\
        );

    \I__3453\ : Odrv12
    port map (
            O => \N__15917\,
            I => \VALID_c\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__15914\,
            I => \VALID_c\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__15911\,
            I => \VALID_c\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__15904\,
            I => \bluejay_data_inst.n14_cascade_\
        );

    \I__3449\ : InMux
    port map (
            O => \N__15901\,
            I => \N__15898\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__15898\,
            I => \N__15895\
        );

    \I__3447\ : Span4Mux_h
    port map (
            O => \N__15895\,
            I => \N__15892\
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__15892\,
            I => n5546
        );

    \I__3445\ : CascadeMux
    port map (
            O => \N__15889\,
            I => \bluejay_data_inst.valid_o_N_155_cascade_\
        );

    \I__3444\ : InMux
    port map (
            O => \N__15886\,
            I => \N__15883\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__15883\,
            I => \bluejay_data_inst.n10\
        );

    \I__3442\ : CascadeMux
    port map (
            O => \N__15880\,
            I => \bluejay_data_inst.n31_cascade_\
        );

    \I__3441\ : CascadeMux
    port map (
            O => \N__15877\,
            I => \bluejay_data_inst.n4253_cascade_\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__15874\,
            I => \bluejay_data_inst.n1038_cascade_\
        );

    \I__3439\ : InMux
    port map (
            O => \N__15871\,
            I => \N__15867\
        );

    \I__3438\ : InMux
    port map (
            O => \N__15870\,
            I => \N__15864\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__15867\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_2\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__15864\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_2\
        );

    \I__3435\ : InMux
    port map (
            O => \N__15859\,
            I => \N__15855\
        );

    \I__3434\ : InMux
    port map (
            O => \N__15858\,
            I => \N__15852\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__15855\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_1\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__15852\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_1\
        );

    \I__3431\ : InMux
    port map (
            O => \N__15847\,
            I => \N__15843\
        );

    \I__3430\ : InMux
    port map (
            O => \N__15846\,
            I => \N__15840\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__15843\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_4\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__15840\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_4\
        );

    \I__3427\ : InMux
    port map (
            O => \N__15835\,
            I => \N__15831\
        );

    \I__3426\ : InMux
    port map (
            O => \N__15834\,
            I => \N__15828\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__15831\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_0\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__15828\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_0\
        );

    \I__3423\ : CascadeMux
    port map (
            O => \N__15823\,
            I => \usb_to_bluejay_if_inst.n12_cascade_\
        );

    \I__3422\ : InMux
    port map (
            O => \N__15820\,
            I => \N__15817\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__15817\,
            I => \usb_to_bluejay_if_inst.n13\
        );

    \I__3420\ : InMux
    port map (
            O => \N__15814\,
            I => \N__15807\
        );

    \I__3419\ : InMux
    port map (
            O => \N__15813\,
            I => \N__15804\
        );

    \I__3418\ : InMux
    port map (
            O => \N__15812\,
            I => \N__15797\
        );

    \I__3417\ : InMux
    port map (
            O => \N__15811\,
            I => \N__15797\
        );

    \I__3416\ : InMux
    port map (
            O => \N__15810\,
            I => \N__15797\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__15807\,
            I => n11
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__15804\,
            I => n11
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__15797\,
            I => n11
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__15790\,
            I => \n11_cascade_\
        );

    \I__3411\ : InMux
    port map (
            O => \N__15787\,
            I => \N__15772\
        );

    \I__3410\ : InMux
    port map (
            O => \N__15786\,
            I => \N__15772\
        );

    \I__3409\ : InMux
    port map (
            O => \N__15785\,
            I => \N__15772\
        );

    \I__3408\ : InMux
    port map (
            O => \N__15784\,
            I => \N__15772\
        );

    \I__3407\ : InMux
    port map (
            O => \N__15783\,
            I => \N__15762\
        );

    \I__3406\ : InMux
    port map (
            O => \N__15782\,
            I => \N__15762\
        );

    \I__3405\ : InMux
    port map (
            O => \N__15781\,
            I => \N__15762\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__15772\,
            I => \N__15759\
        );

    \I__3403\ : InMux
    port map (
            O => \N__15771\,
            I => \N__15750\
        );

    \I__3402\ : InMux
    port map (
            O => \N__15770\,
            I => \N__15745\
        );

    \I__3401\ : InMux
    port map (
            O => \N__15769\,
            I => \N__15745\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__15762\,
            I => \N__15742\
        );

    \I__3399\ : Span4Mux_h
    port map (
            O => \N__15759\,
            I => \N__15739\
        );

    \I__3398\ : InMux
    port map (
            O => \N__15758\,
            I => \N__15734\
        );

    \I__3397\ : InMux
    port map (
            O => \N__15757\,
            I => \N__15734\
        );

    \I__3396\ : InMux
    port map (
            O => \N__15756\,
            I => \N__15725\
        );

    \I__3395\ : InMux
    port map (
            O => \N__15755\,
            I => \N__15725\
        );

    \I__3394\ : InMux
    port map (
            O => \N__15754\,
            I => \N__15725\
        );

    \I__3393\ : InMux
    port map (
            O => \N__15753\,
            I => \N__15725\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__15750\,
            I => state_2_adj_657
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__15745\,
            I => state_2_adj_657
        );

    \I__3390\ : Odrv4
    port map (
            O => \N__15742\,
            I => state_2_adj_657
        );

    \I__3389\ : Odrv4
    port map (
            O => \N__15739\,
            I => state_2_adj_657
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__15734\,
            I => state_2_adj_657
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__15725\,
            I => state_2_adj_657
        );

    \I__3386\ : CascadeMux
    port map (
            O => \N__15712\,
            I => \N__15703\
        );

    \I__3385\ : CascadeMux
    port map (
            O => \N__15711\,
            I => \N__15698\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__15710\,
            I => \N__15695\
        );

    \I__3383\ : InMux
    port map (
            O => \N__15709\,
            I => \N__15692\
        );

    \I__3382\ : InMux
    port map (
            O => \N__15708\,
            I => \N__15686\
        );

    \I__3381\ : InMux
    port map (
            O => \N__15707\,
            I => \N__15686\
        );

    \I__3380\ : InMux
    port map (
            O => \N__15706\,
            I => \N__15677\
        );

    \I__3379\ : InMux
    port map (
            O => \N__15703\,
            I => \N__15670\
        );

    \I__3378\ : InMux
    port map (
            O => \N__15702\,
            I => \N__15670\
        );

    \I__3377\ : InMux
    port map (
            O => \N__15701\,
            I => \N__15670\
        );

    \I__3376\ : InMux
    port map (
            O => \N__15698\,
            I => \N__15667\
        );

    \I__3375\ : InMux
    port map (
            O => \N__15695\,
            I => \N__15664\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__15692\,
            I => \N__15661\
        );

    \I__3373\ : InMux
    port map (
            O => \N__15691\,
            I => \N__15658\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__15686\,
            I => \N__15655\
        );

    \I__3371\ : InMux
    port map (
            O => \N__15685\,
            I => \N__15646\
        );

    \I__3370\ : InMux
    port map (
            O => \N__15684\,
            I => \N__15646\
        );

    \I__3369\ : InMux
    port map (
            O => \N__15683\,
            I => \N__15646\
        );

    \I__3368\ : InMux
    port map (
            O => \N__15682\,
            I => \N__15646\
        );

    \I__3367\ : InMux
    port map (
            O => \N__15681\,
            I => \N__15641\
        );

    \I__3366\ : InMux
    port map (
            O => \N__15680\,
            I => \N__15641\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__15677\,
            I => \N__15636\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__15670\,
            I => \N__15636\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__15667\,
            I => state_1
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__15664\,
            I => state_1
        );

    \I__3361\ : Odrv4
    port map (
            O => \N__15661\,
            I => state_1
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__15658\,
            I => state_1
        );

    \I__3359\ : Odrv4
    port map (
            O => \N__15655\,
            I => state_1
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__15646\,
            I => state_1
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__15641\,
            I => state_1
        );

    \I__3356\ : Odrv4
    port map (
            O => \N__15636\,
            I => state_1
        );

    \I__3355\ : CascadeMux
    port map (
            O => \N__15619\,
            I => \usb_to_bluejay_if_inst.n82_adj_628_cascade_\
        );

    \I__3354\ : InMux
    port map (
            O => \N__15616\,
            I => \N__15609\
        );

    \I__3353\ : InMux
    port map (
            O => \N__15615\,
            I => \N__15609\
        );

    \I__3352\ : InMux
    port map (
            O => \N__15614\,
            I => \N__15606\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__15609\,
            I => \N__15601\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__15606\,
            I => \N__15601\
        );

    \I__3349\ : Odrv4
    port map (
            O => \N__15601\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_7__N_178\
        );

    \I__3348\ : InMux
    port map (
            O => \N__15598\,
            I => \N__15592\
        );

    \I__3347\ : InMux
    port map (
            O => \N__15597\,
            I => \N__15592\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__15592\,
            I => \usb_to_bluejay_if_inst.n2561\
        );

    \I__3345\ : InMux
    port map (
            O => \N__15589\,
            I => \N__15586\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__15586\,
            I => \N__15582\
        );

    \I__3343\ : InMux
    port map (
            O => \N__15585\,
            I => \N__15573\
        );

    \I__3342\ : Span4Mux_h
    port map (
            O => \N__15582\,
            I => \N__15570\
        );

    \I__3341\ : InMux
    port map (
            O => \N__15581\,
            I => \N__15567\
        );

    \I__3340\ : InMux
    port map (
            O => \N__15580\,
            I => \N__15560\
        );

    \I__3339\ : InMux
    port map (
            O => \N__15579\,
            I => \N__15560\
        );

    \I__3338\ : InMux
    port map (
            O => \N__15578\,
            I => \N__15560\
        );

    \I__3337\ : InMux
    port map (
            O => \N__15577\,
            I => \N__15555\
        );

    \I__3336\ : InMux
    port map (
            O => \N__15576\,
            I => \N__15555\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__15573\,
            I => \pc_tx.r_SM_Main_0\
        );

    \I__3334\ : Odrv4
    port map (
            O => \N__15570\,
            I => \pc_tx.r_SM_Main_0\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__15567\,
            I => \pc_tx.r_SM_Main_0\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__15560\,
            I => \pc_tx.r_SM_Main_0\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__15555\,
            I => \pc_tx.r_SM_Main_0\
        );

    \I__3330\ : CascadeMux
    port map (
            O => \N__15544\,
            I => \N__15541\
        );

    \I__3329\ : InMux
    port map (
            O => \N__15541\,
            I => \N__15537\
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__15540\,
            I => \N__15533\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__15537\,
            I => \N__15530\
        );

    \I__3326\ : InMux
    port map (
            O => \N__15536\,
            I => \N__15527\
        );

    \I__3325\ : InMux
    port map (
            O => \N__15533\,
            I => \N__15519\
        );

    \I__3324\ : Span4Mux_h
    port map (
            O => \N__15530\,
            I => \N__15514\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__15527\,
            I => \N__15511\
        );

    \I__3322\ : InMux
    port map (
            O => \N__15526\,
            I => \N__15506\
        );

    \I__3321\ : InMux
    port map (
            O => \N__15525\,
            I => \N__15506\
        );

    \I__3320\ : CascadeMux
    port map (
            O => \N__15524\,
            I => \N__15502\
        );

    \I__3319\ : InMux
    port map (
            O => \N__15523\,
            I => \N__15499\
        );

    \I__3318\ : InMux
    port map (
            O => \N__15522\,
            I => \N__15496\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__15519\,
            I => \N__15493\
        );

    \I__3316\ : InMux
    port map (
            O => \N__15518\,
            I => \N__15488\
        );

    \I__3315\ : InMux
    port map (
            O => \N__15517\,
            I => \N__15488\
        );

    \I__3314\ : Span4Mux_h
    port map (
            O => \N__15514\,
            I => \N__15481\
        );

    \I__3313\ : Span4Mux_h
    port map (
            O => \N__15511\,
            I => \N__15481\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__15506\,
            I => \N__15481\
        );

    \I__3311\ : InMux
    port map (
            O => \N__15505\,
            I => \N__15476\
        );

    \I__3310\ : InMux
    port map (
            O => \N__15502\,
            I => \N__15476\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__15499\,
            I => \r_SM_Main_1_adj_660\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__15496\,
            I => \r_SM_Main_1_adj_660\
        );

    \I__3307\ : Odrv4
    port map (
            O => \N__15493\,
            I => \r_SM_Main_1_adj_660\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__15488\,
            I => \r_SM_Main_1_adj_660\
        );

    \I__3305\ : Odrv4
    port map (
            O => \N__15481\,
            I => \r_SM_Main_1_adj_660\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__15476\,
            I => \r_SM_Main_1_adj_660\
        );

    \I__3303\ : InMux
    port map (
            O => \N__15463\,
            I => \N__15460\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__15460\,
            I => \N__15456\
        );

    \I__3301\ : InMux
    port map (
            O => \N__15459\,
            I => \N__15449\
        );

    \I__3300\ : Span4Mux_h
    port map (
            O => \N__15456\,
            I => \N__15446\
        );

    \I__3299\ : InMux
    port map (
            O => \N__15455\,
            I => \N__15443\
        );

    \I__3298\ : InMux
    port map (
            O => \N__15454\,
            I => \N__15440\
        );

    \I__3297\ : InMux
    port map (
            O => \N__15453\,
            I => \N__15435\
        );

    \I__3296\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15435\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__15449\,
            I => \pc_tx.r_SM_Main_2_N_322_1\
        );

    \I__3294\ : Odrv4
    port map (
            O => \N__15446\,
            I => \pc_tx.r_SM_Main_2_N_322_1\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__15443\,
            I => \pc_tx.r_SM_Main_2_N_322_1\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__15440\,
            I => \pc_tx.r_SM_Main_2_N_322_1\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__15435\,
            I => \pc_tx.r_SM_Main_2_N_322_1\
        );

    \I__3290\ : InMux
    port map (
            O => \N__15424\,
            I => \N__15421\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__15421\,
            I => \N__15418\
        );

    \I__3288\ : Odrv4
    port map (
            O => \N__15418\,
            I => n10_adj_671
        );

    \I__3287\ : InMux
    port map (
            O => \N__15415\,
            I => \N__15412\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__15412\,
            I => n16_adj_672
        );

    \I__3285\ : CascadeMux
    port map (
            O => \N__15409\,
            I => \N__15395\
        );

    \I__3284\ : InMux
    port map (
            O => \N__15408\,
            I => \N__15385\
        );

    \I__3283\ : InMux
    port map (
            O => \N__15407\,
            I => \N__15382\
        );

    \I__3282\ : InMux
    port map (
            O => \N__15406\,
            I => \N__15379\
        );

    \I__3281\ : InMux
    port map (
            O => \N__15405\,
            I => \N__15376\
        );

    \I__3280\ : InMux
    port map (
            O => \N__15404\,
            I => \N__15373\
        );

    \I__3279\ : InMux
    port map (
            O => \N__15403\,
            I => \N__15370\
        );

    \I__3278\ : InMux
    port map (
            O => \N__15402\,
            I => \N__15361\
        );

    \I__3277\ : InMux
    port map (
            O => \N__15401\,
            I => \N__15361\
        );

    \I__3276\ : InMux
    port map (
            O => \N__15400\,
            I => \N__15361\
        );

    \I__3275\ : InMux
    port map (
            O => \N__15399\,
            I => \N__15361\
        );

    \I__3274\ : InMux
    port map (
            O => \N__15398\,
            I => \N__15354\
        );

    \I__3273\ : InMux
    port map (
            O => \N__15395\,
            I => \N__15354\
        );

    \I__3272\ : InMux
    port map (
            O => \N__15394\,
            I => \N__15354\
        );

    \I__3271\ : InMux
    port map (
            O => \N__15393\,
            I => \N__15341\
        );

    \I__3270\ : InMux
    port map (
            O => \N__15392\,
            I => \N__15341\
        );

    \I__3269\ : InMux
    port map (
            O => \N__15391\,
            I => \N__15341\
        );

    \I__3268\ : InMux
    port map (
            O => \N__15390\,
            I => \N__15341\
        );

    \I__3267\ : InMux
    port map (
            O => \N__15389\,
            I => \N__15341\
        );

    \I__3266\ : InMux
    port map (
            O => \N__15388\,
            I => \N__15341\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__15385\,
            I => state_0_adj_658
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__15382\,
            I => state_0_adj_658
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__15379\,
            I => state_0_adj_658
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__15376\,
            I => state_0_adj_658
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__15373\,
            I => state_0_adj_658
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__15370\,
            I => state_0_adj_658
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__15361\,
            I => state_0_adj_658
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__15354\,
            I => state_0_adj_658
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__15341\,
            I => state_0_adj_658
        );

    \I__3256\ : CEMux
    port map (
            O => \N__15322\,
            I => \N__15319\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__15319\,
            I => n5122
        );

    \I__3254\ : InMux
    port map (
            O => \N__15316\,
            I => \usb_to_bluejay_if_inst.n4801\
        );

    \I__3253\ : InMux
    port map (
            O => \N__15313\,
            I => \N__15310\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__15310\,
            I => \N__15306\
        );

    \I__3251\ : InMux
    port map (
            O => \N__15309\,
            I => \N__15303\
        );

    \I__3250\ : Odrv4
    port map (
            O => \N__15306\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_3\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__15303\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_3\
        );

    \I__3248\ : InMux
    port map (
            O => \N__15298\,
            I => \N__15295\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__15295\,
            I => \N__15292\
        );

    \I__3246\ : Odrv4
    port map (
            O => \N__15292\,
            I => \usb_to_bluejay_if_inst.n82\
        );

    \I__3245\ : InMux
    port map (
            O => \N__15289\,
            I => \usb_to_bluejay_if_inst.n4802\
        );

    \I__3244\ : InMux
    port map (
            O => \N__15286\,
            I => \usb_to_bluejay_if_inst.n4803\
        );

    \I__3243\ : InMux
    port map (
            O => \N__15283\,
            I => \N__15277\
        );

    \I__3242\ : InMux
    port map (
            O => \N__15282\,
            I => \N__15277\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__15277\,
            I => \usb_to_bluejay_if_inst.n81\
        );

    \I__3240\ : InMux
    port map (
            O => \N__15274\,
            I => \N__15271\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__15271\,
            I => \N__15267\
        );

    \I__3238\ : InMux
    port map (
            O => \N__15270\,
            I => \N__15264\
        );

    \I__3237\ : Odrv4
    port map (
            O => \N__15267\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_5\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__15264\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_5\
        );

    \I__3235\ : InMux
    port map (
            O => \N__15259\,
            I => \N__15256\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__15256\,
            I => \N__15253\
        );

    \I__3233\ : Odrv12
    port map (
            O => \N__15253\,
            I => \usb_to_bluejay_if_inst.n83\
        );

    \I__3232\ : InMux
    port map (
            O => \N__15250\,
            I => \usb_to_bluejay_if_inst.n4804\
        );

    \I__3231\ : InMux
    port map (
            O => \N__15247\,
            I => \N__15243\
        );

    \I__3230\ : InMux
    port map (
            O => \N__15246\,
            I => \N__15240\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__15243\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_6\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__15240\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_6\
        );

    \I__3227\ : InMux
    port map (
            O => \N__15235\,
            I => \usb_to_bluejay_if_inst.n4805\
        );

    \I__3226\ : InMux
    port map (
            O => \N__15232\,
            I => \usb_to_bluejay_if_inst.n4806\
        );

    \I__3225\ : CascadeMux
    port map (
            O => \N__15229\,
            I => \N__15225\
        );

    \I__3224\ : InMux
    port map (
            O => \N__15228\,
            I => \N__15222\
        );

    \I__3223\ : InMux
    port map (
            O => \N__15225\,
            I => \N__15219\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__15222\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_7\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__15219\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_7\
        );

    \I__3220\ : CEMux
    port map (
            O => \N__15214\,
            I => \N__15210\
        );

    \I__3219\ : CEMux
    port map (
            O => \N__15213\,
            I => \N__15207\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__15210\,
            I => \N__15204\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__15207\,
            I => \N__15201\
        );

    \I__3216\ : Odrv4
    port map (
            O => \N__15204\,
            I => \usb_to_bluejay_if_inst.n2527\
        );

    \I__3215\ : Odrv4
    port map (
            O => \N__15201\,
            I => \usb_to_bluejay_if_inst.n2527\
        );

    \I__3214\ : SRMux
    port map (
            O => \N__15196\,
            I => \N__15193\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__15193\,
            I => \N__15190\
        );

    \I__3212\ : Odrv4
    port map (
            O => \N__15190\,
            I => \usb_to_bluejay_if_inst.n4120\
        );

    \I__3211\ : InMux
    port map (
            O => \N__15187\,
            I => \N__15184\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__15184\,
            I => \N__15181\
        );

    \I__3209\ : Odrv4
    port map (
            O => \N__15181\,
            I => \bluejay_data_inst.n5524\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__15178\,
            I => \N__15175\
        );

    \I__3207\ : InMux
    port map (
            O => \N__15175\,
            I => \N__15172\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__15172\,
            I => \bluejay_data_inst.n1432\
        );

    \I__3205\ : InMux
    port map (
            O => \N__15169\,
            I => \N__15166\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__15166\,
            I => \N__15163\
        );

    \I__3203\ : Span4Mux_v
    port map (
            O => \N__15163\,
            I => \N__15160\
        );

    \I__3202\ : Span4Mux_h
    port map (
            O => \N__15160\,
            I => \N__15157\
        );

    \I__3201\ : Span4Mux_v
    port map (
            O => \N__15157\,
            I => \N__15154\
        );

    \I__3200\ : Sp12to4
    port map (
            O => \N__15154\,
            I => \N__15151\
        );

    \I__3199\ : Odrv12
    port map (
            O => \N__15151\,
            I => \FIFO_D3_c_3\
        );

    \I__3198\ : IoInMux
    port map (
            O => \N__15148\,
            I => \N__15145\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__15145\,
            I => \N__15142\
        );

    \I__3196\ : Span4Mux_s1_v
    port map (
            O => \N__15142\,
            I => \N__15139\
        );

    \I__3195\ : Span4Mux_v
    port map (
            O => \N__15139\,
            I => \N__15136\
        );

    \I__3194\ : Span4Mux_v
    port map (
            O => \N__15136\,
            I => \N__15133\
        );

    \I__3193\ : Span4Mux_v
    port map (
            O => \N__15133\,
            I => \N__15130\
        );

    \I__3192\ : Odrv4
    port map (
            O => \N__15130\,
            I => \DATA3_c_3\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__15127\,
            I => \n3_adj_669_cascade_\
        );

    \I__3190\ : InMux
    port map (
            O => \N__15124\,
            I => \N__15121\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__15121\,
            I => \N__15118\
        );

    \I__3188\ : Span12Mux_v
    port map (
            O => \N__15118\,
            I => \N__15115\
        );

    \I__3187\ : Span12Mux_h
    port map (
            O => \N__15115\,
            I => \N__15112\
        );

    \I__3186\ : Odrv12
    port map (
            O => \N__15112\,
            I => \FIFO_D12_c_12\
        );

    \I__3185\ : IoInMux
    port map (
            O => \N__15109\,
            I => \N__15106\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__15106\,
            I => \N__15103\
        );

    \I__3183\ : Span4Mux_s2_h
    port map (
            O => \N__15103\,
            I => \N__15100\
        );

    \I__3182\ : Span4Mux_v
    port map (
            O => \N__15100\,
            I => \N__15097\
        );

    \I__3181\ : Sp12to4
    port map (
            O => \N__15097\,
            I => \N__15094\
        );

    \I__3180\ : Odrv12
    port map (
            O => \N__15094\,
            I => \DATA12_c_12\
        );

    \I__3179\ : InMux
    port map (
            O => \N__15091\,
            I => \N__15080\
        );

    \I__3178\ : InMux
    port map (
            O => \N__15090\,
            I => \N__15071\
        );

    \I__3177\ : InMux
    port map (
            O => \N__15089\,
            I => \N__15071\
        );

    \I__3176\ : InMux
    port map (
            O => \N__15088\,
            I => \N__15071\
        );

    \I__3175\ : InMux
    port map (
            O => \N__15087\,
            I => \N__15071\
        );

    \I__3174\ : InMux
    port map (
            O => \N__15086\,
            I => \N__15068\
        );

    \I__3173\ : InMux
    port map (
            O => \N__15085\,
            I => \N__15061\
        );

    \I__3172\ : InMux
    port map (
            O => \N__15084\,
            I => \N__15061\
        );

    \I__3171\ : InMux
    port map (
            O => \N__15083\,
            I => \N__15061\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__15080\,
            I => \N__15055\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__15071\,
            I => \N__15048\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__15068\,
            I => \N__15043\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__15061\,
            I => \N__15043\
        );

    \I__3166\ : InMux
    port map (
            O => \N__15060\,
            I => \N__15036\
        );

    \I__3165\ : InMux
    port map (
            O => \N__15059\,
            I => \N__15036\
        );

    \I__3164\ : InMux
    port map (
            O => \N__15058\,
            I => \N__15036\
        );

    \I__3163\ : Span4Mux_v
    port map (
            O => \N__15055\,
            I => \N__15033\
        );

    \I__3162\ : InMux
    port map (
            O => \N__15054\,
            I => \N__15030\
        );

    \I__3161\ : InMux
    port map (
            O => \N__15053\,
            I => \N__15023\
        );

    \I__3160\ : InMux
    port map (
            O => \N__15052\,
            I => \N__15023\
        );

    \I__3159\ : InMux
    port map (
            O => \N__15051\,
            I => \N__15023\
        );

    \I__3158\ : Span4Mux_h
    port map (
            O => \N__15048\,
            I => \N__15018\
        );

    \I__3157\ : Span4Mux_h
    port map (
            O => \N__15043\,
            I => \N__15013\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__15036\,
            I => \N__15013\
        );

    \I__3155\ : Sp12to4
    port map (
            O => \N__15033\,
            I => \N__15006\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__15030\,
            I => \N__15006\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__15023\,
            I => \N__15006\
        );

    \I__3152\ : InMux
    port map (
            O => \N__15022\,
            I => \N__15003\
        );

    \I__3151\ : InMux
    port map (
            O => \N__15021\,
            I => \N__15000\
        );

    \I__3150\ : Odrv4
    port map (
            O => \N__15018\,
            I => uart_rx_complete_rising_edge
        );

    \I__3149\ : Odrv4
    port map (
            O => \N__15013\,
            I => uart_rx_complete_rising_edge
        );

    \I__3148\ : Odrv12
    port map (
            O => \N__15006\,
            I => uart_rx_complete_rising_edge
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__15003\,
            I => uart_rx_complete_rising_edge
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__15000\,
            I => uart_rx_complete_rising_edge
        );

    \I__3145\ : InMux
    port map (
            O => \N__14989\,
            I => \N__14985\
        );

    \I__3144\ : InMux
    port map (
            O => \N__14988\,
            I => \N__14982\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__14985\,
            I => even_byte_flag
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__14982\,
            I => even_byte_flag
        );

    \I__3141\ : InMux
    port map (
            O => \N__14977\,
            I => \bfn_16_5_0_\
        );

    \I__3140\ : InMux
    port map (
            O => \N__14974\,
            I => \usb_to_bluejay_if_inst.n4800\
        );

    \I__3139\ : CascadeMux
    port map (
            O => \N__14971\,
            I => \N__14966\
        );

    \I__3138\ : InMux
    port map (
            O => \N__14970\,
            I => \N__14963\
        );

    \I__3137\ : InMux
    port map (
            O => \N__14969\,
            I => \N__14960\
        );

    \I__3136\ : InMux
    port map (
            O => \N__14966\,
            I => \N__14957\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__14963\,
            I => \bluejay_data_inst.v_counter_9\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__14960\,
            I => \bluejay_data_inst.v_counter_9\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__14957\,
            I => \bluejay_data_inst.v_counter_9\
        );

    \I__3132\ : InMux
    port map (
            O => \N__14950\,
            I => \N__14947\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__14947\,
            I => \bluejay_data_inst.n1100\
        );

    \I__3130\ : InMux
    port map (
            O => \N__14944\,
            I => \bluejay_data_inst.n4856\
        );

    \I__3129\ : InMux
    port map (
            O => \N__14941\,
            I => \N__14936\
        );

    \I__3128\ : InMux
    port map (
            O => \N__14940\,
            I => \N__14933\
        );

    \I__3127\ : InMux
    port map (
            O => \N__14939\,
            I => \N__14930\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__14936\,
            I => \bluejay_data_inst.v_counter_10\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__14933\,
            I => \bluejay_data_inst.v_counter_10\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__14930\,
            I => \bluejay_data_inst.v_counter_10\
        );

    \I__3123\ : InMux
    port map (
            O => \N__14923\,
            I => \bluejay_data_inst.n4857\
        );

    \I__3122\ : InMux
    port map (
            O => \N__14920\,
            I => \N__14917\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__14917\,
            I => \bluejay_data_inst.n1099\
        );

    \I__3120\ : CascadeMux
    port map (
            O => \N__14914\,
            I => \bluejay_data_inst.n1054_cascade_\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__14911\,
            I => \N__14904\
        );

    \I__3118\ : CascadeMux
    port map (
            O => \N__14910\,
            I => \N__14901\
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__14909\,
            I => \N__14898\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__14908\,
            I => \N__14891\
        );

    \I__3115\ : CascadeMux
    port map (
            O => \N__14907\,
            I => \N__14887\
        );

    \I__3114\ : InMux
    port map (
            O => \N__14904\,
            I => \N__14880\
        );

    \I__3113\ : InMux
    port map (
            O => \N__14901\,
            I => \N__14880\
        );

    \I__3112\ : InMux
    port map (
            O => \N__14898\,
            I => \N__14880\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__14897\,
            I => \N__14877\
        );

    \I__3110\ : CascadeMux
    port map (
            O => \N__14896\,
            I => \N__14873\
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__14895\,
            I => \N__14870\
        );

    \I__3108\ : InMux
    port map (
            O => \N__14894\,
            I => \N__14866\
        );

    \I__3107\ : InMux
    port map (
            O => \N__14891\,
            I => \N__14859\
        );

    \I__3106\ : InMux
    port map (
            O => \N__14890\,
            I => \N__14859\
        );

    \I__3105\ : InMux
    port map (
            O => \N__14887\,
            I => \N__14859\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__14880\,
            I => \N__14856\
        );

    \I__3103\ : InMux
    port map (
            O => \N__14877\,
            I => \N__14845\
        );

    \I__3102\ : InMux
    port map (
            O => \N__14876\,
            I => \N__14845\
        );

    \I__3101\ : InMux
    port map (
            O => \N__14873\,
            I => \N__14845\
        );

    \I__3100\ : InMux
    port map (
            O => \N__14870\,
            I => \N__14845\
        );

    \I__3099\ : InMux
    port map (
            O => \N__14869\,
            I => \N__14845\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__14866\,
            I => \bluejay_data_inst.n1373\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__14859\,
            I => \bluejay_data_inst.n1373\
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__14856\,
            I => \bluejay_data_inst.n1373\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__14845\,
            I => \bluejay_data_inst.n1373\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__14836\,
            I => \n5_cascade_\
        );

    \I__3093\ : InMux
    port map (
            O => \N__14833\,
            I => \N__14828\
        );

    \I__3092\ : InMux
    port map (
            O => \N__14832\,
            I => \N__14825\
        );

    \I__3091\ : InMux
    port map (
            O => \N__14831\,
            I => \N__14822\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__14828\,
            I => \bluejay_data_inst.v_counter_1\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__14825\,
            I => \bluejay_data_inst.v_counter_1\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__14822\,
            I => \bluejay_data_inst.v_counter_1\
        );

    \I__3087\ : InMux
    port map (
            O => \N__14815\,
            I => \N__14812\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__14812\,
            I => \bluejay_data_inst.n1108\
        );

    \I__3085\ : InMux
    port map (
            O => \N__14809\,
            I => \bluejay_data_inst.n4848\
        );

    \I__3084\ : InMux
    port map (
            O => \N__14806\,
            I => \N__14801\
        );

    \I__3083\ : InMux
    port map (
            O => \N__14805\,
            I => \N__14798\
        );

    \I__3082\ : InMux
    port map (
            O => \N__14804\,
            I => \N__14795\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__14801\,
            I => \bluejay_data_inst.v_counter_2\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__14798\,
            I => \bluejay_data_inst.v_counter_2\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__14795\,
            I => \bluejay_data_inst.v_counter_2\
        );

    \I__3078\ : InMux
    port map (
            O => \N__14788\,
            I => \N__14785\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__14785\,
            I => \bluejay_data_inst.n1107\
        );

    \I__3076\ : InMux
    port map (
            O => \N__14782\,
            I => \bluejay_data_inst.n4849\
        );

    \I__3075\ : InMux
    port map (
            O => \N__14779\,
            I => \N__14774\
        );

    \I__3074\ : InMux
    port map (
            O => \N__14778\,
            I => \N__14771\
        );

    \I__3073\ : InMux
    port map (
            O => \N__14777\,
            I => \N__14768\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__14774\,
            I => \bluejay_data_inst.v_counter_3\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__14771\,
            I => \bluejay_data_inst.v_counter_3\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__14768\,
            I => \bluejay_data_inst.v_counter_3\
        );

    \I__3069\ : InMux
    port map (
            O => \N__14761\,
            I => \N__14758\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__14758\,
            I => \bluejay_data_inst.n1106\
        );

    \I__3067\ : InMux
    port map (
            O => \N__14755\,
            I => \bluejay_data_inst.n4850\
        );

    \I__3066\ : InMux
    port map (
            O => \N__14752\,
            I => \N__14749\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__14749\,
            I => \N__14746\
        );

    \I__3064\ : Span4Mux_h
    port map (
            O => \N__14746\,
            I => \N__14741\
        );

    \I__3063\ : InMux
    port map (
            O => \N__14745\,
            I => \N__14736\
        );

    \I__3062\ : InMux
    port map (
            O => \N__14744\,
            I => \N__14736\
        );

    \I__3061\ : Odrv4
    port map (
            O => \N__14741\,
            I => \bluejay_data_inst.v_counter_4\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__14736\,
            I => \bluejay_data_inst.v_counter_4\
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__14731\,
            I => \N__14728\
        );

    \I__3058\ : InMux
    port map (
            O => \N__14728\,
            I => \N__14725\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__14725\,
            I => \N__14722\
        );

    \I__3056\ : Odrv4
    port map (
            O => \N__14722\,
            I => \bluejay_data_inst.n1105\
        );

    \I__3055\ : InMux
    port map (
            O => \N__14719\,
            I => \bluejay_data_inst.n4851\
        );

    \I__3054\ : CascadeMux
    port map (
            O => \N__14716\,
            I => \N__14713\
        );

    \I__3053\ : InMux
    port map (
            O => \N__14713\,
            I => \N__14709\
        );

    \I__3052\ : CascadeMux
    port map (
            O => \N__14712\,
            I => \N__14705\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__14709\,
            I => \N__14702\
        );

    \I__3050\ : InMux
    port map (
            O => \N__14708\,
            I => \N__14697\
        );

    \I__3049\ : InMux
    port map (
            O => \N__14705\,
            I => \N__14697\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__14702\,
            I => \bluejay_data_inst.v_counter_5\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__14697\,
            I => \bluejay_data_inst.v_counter_5\
        );

    \I__3046\ : InMux
    port map (
            O => \N__14692\,
            I => \N__14689\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__14689\,
            I => \N__14686\
        );

    \I__3044\ : Odrv4
    port map (
            O => \N__14686\,
            I => \bluejay_data_inst.n1104\
        );

    \I__3043\ : InMux
    port map (
            O => \N__14683\,
            I => \bluejay_data_inst.n4852\
        );

    \I__3042\ : InMux
    port map (
            O => \N__14680\,
            I => \N__14675\
        );

    \I__3041\ : InMux
    port map (
            O => \N__14679\,
            I => \N__14672\
        );

    \I__3040\ : InMux
    port map (
            O => \N__14678\,
            I => \N__14669\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__14675\,
            I => \bluejay_data_inst.v_counter_6\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__14672\,
            I => \bluejay_data_inst.v_counter_6\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__14669\,
            I => \bluejay_data_inst.v_counter_6\
        );

    \I__3036\ : InMux
    port map (
            O => \N__14662\,
            I => \N__14659\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__14659\,
            I => \bluejay_data_inst.n1103\
        );

    \I__3034\ : InMux
    port map (
            O => \N__14656\,
            I => \bluejay_data_inst.n4853\
        );

    \I__3033\ : InMux
    port map (
            O => \N__14653\,
            I => \N__14650\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__14650\,
            I => \N__14645\
        );

    \I__3031\ : InMux
    port map (
            O => \N__14649\,
            I => \N__14642\
        );

    \I__3030\ : InMux
    port map (
            O => \N__14648\,
            I => \N__14639\
        );

    \I__3029\ : Odrv4
    port map (
            O => \N__14645\,
            I => \bluejay_data_inst.v_counter_7\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__14642\,
            I => \bluejay_data_inst.v_counter_7\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__14639\,
            I => \bluejay_data_inst.v_counter_7\
        );

    \I__3026\ : InMux
    port map (
            O => \N__14632\,
            I => \N__14629\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__14629\,
            I => \bluejay_data_inst.n1102\
        );

    \I__3024\ : InMux
    port map (
            O => \N__14626\,
            I => \bfn_15_9_0_\
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__14623\,
            I => \N__14619\
        );

    \I__3022\ : InMux
    port map (
            O => \N__14622\,
            I => \N__14615\
        );

    \I__3021\ : InMux
    port map (
            O => \N__14619\,
            I => \N__14612\
        );

    \I__3020\ : InMux
    port map (
            O => \N__14618\,
            I => \N__14609\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__14615\,
            I => \bluejay_data_inst.v_counter_8\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__14612\,
            I => \bluejay_data_inst.v_counter_8\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__14609\,
            I => \bluejay_data_inst.v_counter_8\
        );

    \I__3016\ : InMux
    port map (
            O => \N__14602\,
            I => \N__14599\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__14599\,
            I => \bluejay_data_inst.n1101\
        );

    \I__3014\ : InMux
    port map (
            O => \N__14596\,
            I => \bluejay_data_inst.n4855\
        );

    \I__3013\ : CascadeMux
    port map (
            O => \N__14593\,
            I => \usb_to_bluejay_if_inst.n2492_cascade_\
        );

    \I__3012\ : CEMux
    port map (
            O => \N__14590\,
            I => \N__14587\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__14587\,
            I => \N__14584\
        );

    \I__3010\ : Odrv4
    port map (
            O => \N__14584\,
            I => \usb_to_bluejay_if_inst.n2492\
        );

    \I__3009\ : SRMux
    port map (
            O => \N__14581\,
            I => \N__14578\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__14578\,
            I => \N__14575\
        );

    \I__3007\ : Odrv4
    port map (
            O => \N__14575\,
            I => \usb_to_bluejay_if_inst.n4963\
        );

    \I__3006\ : InMux
    port map (
            O => \N__14572\,
            I => \N__14564\
        );

    \I__3005\ : InMux
    port map (
            O => \N__14571\,
            I => \N__14564\
        );

    \I__3004\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14560\
        );

    \I__3003\ : InMux
    port map (
            O => \N__14569\,
            I => \N__14557\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__14564\,
            I => \N__14554\
        );

    \I__3001\ : InMux
    port map (
            O => \N__14563\,
            I => \N__14551\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__14560\,
            I => \usb_to_bluejay_if_inst.n3\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__14557\,
            I => \usb_to_bluejay_if_inst.n3\
        );

    \I__2998\ : Odrv4
    port map (
            O => \N__14554\,
            I => \usb_to_bluejay_if_inst.n3\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__14551\,
            I => \usb_to_bluejay_if_inst.n3\
        );

    \I__2996\ : CascadeMux
    port map (
            O => \N__14542\,
            I => \usb_to_bluejay_if_inst.state_timeout_counter_7__N_178_cascade_\
        );

    \I__2995\ : InMux
    port map (
            O => \N__14539\,
            I => \N__14536\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__14536\,
            I => \usb_to_bluejay_if_inst.n5400\
        );

    \I__2993\ : CascadeMux
    port map (
            O => \N__14533\,
            I => \usb_to_bluejay_if_inst.n2562_cascade_\
        );

    \I__2992\ : InMux
    port map (
            O => \N__14530\,
            I => \N__14527\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__14527\,
            I => \usb_to_bluejay_if_inst.n2564\
        );

    \I__2990\ : CascadeMux
    port map (
            O => \N__14524\,
            I => \usb_to_bluejay_if_inst.n2564_cascade_\
        );

    \I__2989\ : SRMux
    port map (
            O => \N__14521\,
            I => \N__14518\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__14518\,
            I => \N__14515\
        );

    \I__2987\ : Odrv12
    port map (
            O => \N__14515\,
            I => \usb_to_bluejay_if_inst.n2706\
        );

    \I__2986\ : InMux
    port map (
            O => \N__14512\,
            I => \N__14507\
        );

    \I__2985\ : InMux
    port map (
            O => \N__14511\,
            I => \N__14504\
        );

    \I__2984\ : InMux
    port map (
            O => \N__14510\,
            I => \N__14501\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__14507\,
            I => \bluejay_data_inst.v_counter_0\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__14504\,
            I => \bluejay_data_inst.v_counter_0\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__14501\,
            I => \bluejay_data_inst.v_counter_0\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__14494\,
            I => \N__14491\
        );

    \I__2979\ : InMux
    port map (
            O => \N__14491\,
            I => \N__14488\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__14488\,
            I => \bluejay_data_inst.n1476\
        );

    \I__2977\ : InMux
    port map (
            O => \N__14485\,
            I => \N__14482\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__14482\,
            I => \bluejay_data_inst.n1109\
        );

    \I__2975\ : InMux
    port map (
            O => \N__14479\,
            I => \bluejay_data_inst.n4847\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__14476\,
            I => \N__14472\
        );

    \I__2973\ : InMux
    port map (
            O => \N__14475\,
            I => \N__14469\
        );

    \I__2972\ : InMux
    port map (
            O => \N__14472\,
            I => \N__14466\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__14469\,
            I => \N__14463\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__14466\,
            I => \N__14460\
        );

    \I__2969\ : Span4Mux_h
    port map (
            O => \N__14463\,
            I => \N__14457\
        );

    \I__2968\ : Span4Mux_h
    port map (
            O => \N__14460\,
            I => \N__14454\
        );

    \I__2967\ : Span4Mux_v
    port map (
            O => \N__14457\,
            I => \N__14449\
        );

    \I__2966\ : Span4Mux_h
    port map (
            O => \N__14454\,
            I => \N__14449\
        );

    \I__2965\ : Odrv4
    port map (
            O => \N__14449\,
            I => n5_adj_667
        );

    \I__2964\ : InMux
    port map (
            O => \N__14446\,
            I => \N__14443\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__14443\,
            I => \N__14440\
        );

    \I__2962\ : Span4Mux_v
    port map (
            O => \N__14440\,
            I => \N__14437\
        );

    \I__2961\ : Span4Mux_h
    port map (
            O => \N__14437\,
            I => \N__14433\
        );

    \I__2960\ : InMux
    port map (
            O => \N__14436\,
            I => \N__14430\
        );

    \I__2959\ : Odrv4
    port map (
            O => \N__14433\,
            I => start_transfer_edge
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__14430\,
            I => start_transfer_edge
        );

    \I__2957\ : CascadeMux
    port map (
            O => \N__14425\,
            I => \usb_to_bluejay_if_inst.n5400_cascade_\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__14422\,
            I => \usb_to_bluejay_if_inst.n2527_cascade_\
        );

    \I__2955\ : InMux
    port map (
            O => \N__14419\,
            I => \N__14413\
        );

    \I__2954\ : InMux
    port map (
            O => \N__14418\,
            I => \N__14413\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__14413\,
            I => \N__14410\
        );

    \I__2952\ : Odrv4
    port map (
            O => \N__14410\,
            I => spi_start_transfer_r
        );

    \I__2951\ : InMux
    port map (
            O => \N__14407\,
            I => \N__14404\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__14404\,
            I => start_transfer_prev
        );

    \I__2949\ : InMux
    port map (
            O => \N__14401\,
            I => \N__14396\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__14400\,
            I => \N__14393\
        );

    \I__2947\ : InMux
    port map (
            O => \N__14399\,
            I => \N__14389\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__14396\,
            I => \N__14386\
        );

    \I__2945\ : InMux
    port map (
            O => \N__14393\,
            I => \N__14383\
        );

    \I__2944\ : InMux
    port map (
            O => \N__14392\,
            I => \N__14380\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__14389\,
            I => data_in_fifo_prev
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__14386\,
            I => data_in_fifo_prev
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__14383\,
            I => data_in_fifo_prev
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__14380\,
            I => data_in_fifo_prev
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__14371\,
            I => \usb_to_bluejay_if_inst.n4136_cascade_\
        );

    \I__2938\ : InMux
    port map (
            O => \N__14368\,
            I => \N__14365\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__14365\,
            I => \N__14359\
        );

    \I__2936\ : InMux
    port map (
            O => \N__14364\,
            I => \N__14354\
        );

    \I__2935\ : InMux
    port map (
            O => \N__14363\,
            I => \N__14354\
        );

    \I__2934\ : InMux
    port map (
            O => \N__14362\,
            I => \N__14348\
        );

    \I__2933\ : Span4Mux_h
    port map (
            O => \N__14359\,
            I => \N__14345\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__14354\,
            I => \N__14342\
        );

    \I__2931\ : InMux
    port map (
            O => \N__14353\,
            I => \N__14339\
        );

    \I__2930\ : InMux
    port map (
            O => \N__14352\,
            I => \N__14336\
        );

    \I__2929\ : InMux
    port map (
            O => \N__14351\,
            I => \N__14333\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__14348\,
            I => fifo_read_cmd
        );

    \I__2927\ : Odrv4
    port map (
            O => \N__14345\,
            I => fifo_read_cmd
        );

    \I__2926\ : Odrv4
    port map (
            O => \N__14342\,
            I => fifo_read_cmd
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__14339\,
            I => fifo_read_cmd
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__14336\,
            I => fifo_read_cmd
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__14333\,
            I => fifo_read_cmd
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__14320\,
            I => \N__14315\
        );

    \I__2921\ : InMux
    port map (
            O => \N__14319\,
            I => \N__14312\
        );

    \I__2920\ : InMux
    port map (
            O => \N__14318\,
            I => \N__14309\
        );

    \I__2919\ : InMux
    port map (
            O => \N__14315\,
            I => \N__14306\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__14312\,
            I => \N__14303\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__14309\,
            I => \N__14293\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__14306\,
            I => \N__14293\
        );

    \I__2915\ : Span4Mux_h
    port map (
            O => \N__14303\,
            I => \N__14290\
        );

    \I__2914\ : InMux
    port map (
            O => \N__14302\,
            I => \N__14285\
        );

    \I__2913\ : InMux
    port map (
            O => \N__14301\,
            I => \N__14285\
        );

    \I__2912\ : InMux
    port map (
            O => \N__14300\,
            I => \N__14280\
        );

    \I__2911\ : InMux
    port map (
            O => \N__14299\,
            I => \N__14280\
        );

    \I__2910\ : InMux
    port map (
            O => \N__14298\,
            I => \N__14277\
        );

    \I__2909\ : Odrv12
    port map (
            O => \N__14293\,
            I => is_fifo_empty_flag
        );

    \I__2908\ : Odrv4
    port map (
            O => \N__14290\,
            I => is_fifo_empty_flag
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__14285\,
            I => is_fifo_empty_flag
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__14280\,
            I => is_fifo_empty_flag
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__14277\,
            I => is_fifo_empty_flag
        );

    \I__2904\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14262\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__14265\,
            I => \N__14254\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__14262\,
            I => \N__14251\
        );

    \I__2901\ : InMux
    port map (
            O => \N__14261\,
            I => \N__14248\
        );

    \I__2900\ : InMux
    port map (
            O => \N__14260\,
            I => \N__14243\
        );

    \I__2899\ : InMux
    port map (
            O => \N__14259\,
            I => \N__14240\
        );

    \I__2898\ : InMux
    port map (
            O => \N__14258\,
            I => \N__14237\
        );

    \I__2897\ : InMux
    port map (
            O => \N__14257\,
            I => \N__14234\
        );

    \I__2896\ : InMux
    port map (
            O => \N__14254\,
            I => \N__14230\
        );

    \I__2895\ : Span4Mux_v
    port map (
            O => \N__14251\,
            I => \N__14225\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__14248\,
            I => \N__14225\
        );

    \I__2893\ : CascadeMux
    port map (
            O => \N__14247\,
            I => \N__14222\
        );

    \I__2892\ : InMux
    port map (
            O => \N__14246\,
            I => \N__14218\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__14243\,
            I => \N__14209\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__14240\,
            I => \N__14209\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__14237\,
            I => \N__14209\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__14234\,
            I => \N__14209\
        );

    \I__2887\ : InMux
    port map (
            O => \N__14233\,
            I => \N__14205\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__14230\,
            I => \N__14200\
        );

    \I__2885\ : Span4Mux_h
    port map (
            O => \N__14225\,
            I => \N__14200\
        );

    \I__2884\ : InMux
    port map (
            O => \N__14222\,
            I => \N__14193\
        );

    \I__2883\ : InMux
    port map (
            O => \N__14221\,
            I => \N__14193\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__14218\,
            I => \N__14190\
        );

    \I__2881\ : Span4Mux_v
    port map (
            O => \N__14209\,
            I => \N__14187\
        );

    \I__2880\ : InMux
    port map (
            O => \N__14208\,
            I => \N__14184\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__14205\,
            I => \N__14179\
        );

    \I__2878\ : Span4Mux_v
    port map (
            O => \N__14200\,
            I => \N__14179\
        );

    \I__2877\ : InMux
    port map (
            O => \N__14199\,
            I => \N__14176\
        );

    \I__2876\ : InMux
    port map (
            O => \N__14198\,
            I => \N__14173\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__14193\,
            I => \N__14164\
        );

    \I__2874\ : Span4Mux_v
    port map (
            O => \N__14190\,
            I => \N__14164\
        );

    \I__2873\ : Span4Mux_h
    port map (
            O => \N__14187\,
            I => \N__14164\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__14184\,
            I => \N__14164\
        );

    \I__2871\ : Span4Mux_h
    port map (
            O => \N__14179\,
            I => \N__14161\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__14176\,
            I => \N__14158\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__14173\,
            I => rd_addr_r_0
        );

    \I__2868\ : Odrv4
    port map (
            O => \N__14164\,
            I => rd_addr_r_0
        );

    \I__2867\ : Odrv4
    port map (
            O => \N__14161\,
            I => rd_addr_r_0
        );

    \I__2866\ : Odrv12
    port map (
            O => \N__14158\,
            I => rd_addr_r_0
        );

    \I__2865\ : InMux
    port map (
            O => \N__14149\,
            I => \N__14146\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__14146\,
            I => \N__14143\
        );

    \I__2863\ : Span4Mux_v
    port map (
            O => \N__14143\,
            I => \N__14140\
        );

    \I__2862\ : Sp12to4
    port map (
            O => \N__14140\,
            I => \N__14137\
        );

    \I__2861\ : Span12Mux_h
    port map (
            O => \N__14137\,
            I => \N__14134\
        );

    \I__2860\ : Span12Mux_v
    port map (
            O => \N__14134\,
            I => \N__14131\
        );

    \I__2859\ : Odrv12
    port map (
            O => \N__14131\,
            I => \FIFO_D10_c_10\
        );

    \I__2858\ : IoInMux
    port map (
            O => \N__14128\,
            I => \N__14125\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__14125\,
            I => \N__14122\
        );

    \I__2856\ : IoSpan4Mux
    port map (
            O => \N__14122\,
            I => \N__14119\
        );

    \I__2855\ : Sp12to4
    port map (
            O => \N__14119\,
            I => \N__14116\
        );

    \I__2854\ : Span12Mux_s7_h
    port map (
            O => \N__14116\,
            I => \N__14113\
        );

    \I__2853\ : Odrv12
    port map (
            O => \N__14113\,
            I => \DATA10_c_10\
        );

    \I__2852\ : InMux
    port map (
            O => \N__14110\,
            I => \N__14107\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__14107\,
            I => \N__14104\
        );

    \I__2850\ : Span4Mux_v
    port map (
            O => \N__14104\,
            I => \N__14101\
        );

    \I__2849\ : Sp12to4
    port map (
            O => \N__14101\,
            I => \N__14098\
        );

    \I__2848\ : Span12Mux_h
    port map (
            O => \N__14098\,
            I => \N__14095\
        );

    \I__2847\ : Span12Mux_v
    port map (
            O => \N__14095\,
            I => \N__14092\
        );

    \I__2846\ : Odrv12
    port map (
            O => \N__14092\,
            I => \FIFO_D9_c_9\
        );

    \I__2845\ : IoInMux
    port map (
            O => \N__14089\,
            I => \N__14086\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__14086\,
            I => \N__14083\
        );

    \I__2843\ : IoSpan4Mux
    port map (
            O => \N__14083\,
            I => \N__14080\
        );

    \I__2842\ : IoSpan4Mux
    port map (
            O => \N__14080\,
            I => \N__14077\
        );

    \I__2841\ : Span4Mux_s3_h
    port map (
            O => \N__14077\,
            I => \N__14074\
        );

    \I__2840\ : Sp12to4
    port map (
            O => \N__14074\,
            I => \N__14071\
        );

    \I__2839\ : Odrv12
    port map (
            O => \N__14071\,
            I => \DATA9_c_9\
        );

    \I__2838\ : InMux
    port map (
            O => \N__14068\,
            I => \N__14065\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__14065\,
            I => \N__14062\
        );

    \I__2836\ : Span4Mux_h
    port map (
            O => \N__14062\,
            I => \N__14059\
        );

    \I__2835\ : Sp12to4
    port map (
            O => \N__14059\,
            I => \N__14056\
        );

    \I__2834\ : Span12Mux_v
    port map (
            O => \N__14056\,
            I => \N__14053\
        );

    \I__2833\ : Span12Mux_v
    port map (
            O => \N__14053\,
            I => \N__14050\
        );

    \I__2832\ : Span12Mux_h
    port map (
            O => \N__14050\,
            I => \N__14047\
        );

    \I__2831\ : Odrv12
    port map (
            O => \N__14047\,
            I => \FIFO_D16_c_16\
        );

    \I__2830\ : IoInMux
    port map (
            O => \N__14044\,
            I => \N__14041\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__14041\,
            I => \N__14038\
        );

    \I__2828\ : Span4Mux_s3_h
    port map (
            O => \N__14038\,
            I => \N__14035\
        );

    \I__2827\ : Span4Mux_v
    port map (
            O => \N__14035\,
            I => \N__14032\
        );

    \I__2826\ : Span4Mux_v
    port map (
            O => \N__14032\,
            I => \N__14029\
        );

    \I__2825\ : Sp12to4
    port map (
            O => \N__14029\,
            I => \N__14026\
        );

    \I__2824\ : Odrv12
    port map (
            O => \N__14026\,
            I => \DATA16_c_16\
        );

    \I__2823\ : InMux
    port map (
            O => \N__14023\,
            I => \N__14020\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__14020\,
            I => \N__14013\
        );

    \I__2821\ : InMux
    port map (
            O => \N__14019\,
            I => \N__14010\
        );

    \I__2820\ : InMux
    port map (
            O => \N__14018\,
            I => \N__14006\
        );

    \I__2819\ : InMux
    port map (
            O => \N__14017\,
            I => \N__14003\
        );

    \I__2818\ : InMux
    port map (
            O => \N__14016\,
            I => \N__14000\
        );

    \I__2817\ : Span4Mux_v
    port map (
            O => \N__14013\,
            I => \N__13995\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__14010\,
            I => \N__13995\
        );

    \I__2815\ : InMux
    port map (
            O => \N__14009\,
            I => \N__13992\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__14006\,
            I => \pc_rx.r_Bit_Index_2\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__14003\,
            I => \pc_rx.r_Bit_Index_2\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__14000\,
            I => \pc_rx.r_Bit_Index_2\
        );

    \I__2811\ : Odrv4
    port map (
            O => \N__13995\,
            I => \pc_rx.r_Bit_Index_2\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__13992\,
            I => \pc_rx.r_Bit_Index_2\
        );

    \I__2809\ : InMux
    port map (
            O => \N__13981\,
            I => \N__13969\
        );

    \I__2808\ : InMux
    port map (
            O => \N__13980\,
            I => \N__13969\
        );

    \I__2807\ : InMux
    port map (
            O => \N__13979\,
            I => \N__13964\
        );

    \I__2806\ : InMux
    port map (
            O => \N__13978\,
            I => \N__13964\
        );

    \I__2805\ : InMux
    port map (
            O => \N__13977\,
            I => \N__13961\
        );

    \I__2804\ : InMux
    port map (
            O => \N__13976\,
            I => \N__13956\
        );

    \I__2803\ : InMux
    port map (
            O => \N__13975\,
            I => \N__13956\
        );

    \I__2802\ : InMux
    port map (
            O => \N__13974\,
            I => \N__13953\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__13969\,
            I => \r_Bit_Index_0\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__13964\,
            I => \r_Bit_Index_0\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__13961\,
            I => \r_Bit_Index_0\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__13956\,
            I => \r_Bit_Index_0\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__13953\,
            I => \r_Bit_Index_0\
        );

    \I__2796\ : InMux
    port map (
            O => \N__13942\,
            I => \N__13939\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__13939\,
            I => \N__13931\
        );

    \I__2794\ : InMux
    port map (
            O => \N__13938\,
            I => \N__13928\
        );

    \I__2793\ : InMux
    port map (
            O => \N__13937\,
            I => \N__13922\
        );

    \I__2792\ : InMux
    port map (
            O => \N__13936\,
            I => \N__13922\
        );

    \I__2791\ : InMux
    port map (
            O => \N__13935\,
            I => \N__13917\
        );

    \I__2790\ : InMux
    port map (
            O => \N__13934\,
            I => \N__13917\
        );

    \I__2789\ : Span4Mux_v
    port map (
            O => \N__13931\,
            I => \N__13912\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__13928\,
            I => \N__13912\
        );

    \I__2787\ : InMux
    port map (
            O => \N__13927\,
            I => \N__13909\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__13922\,
            I => \pc_rx.r_Bit_Index_1\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__13917\,
            I => \pc_rx.r_Bit_Index_1\
        );

    \I__2784\ : Odrv4
    port map (
            O => \N__13912\,
            I => \pc_rx.r_Bit_Index_1\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__13909\,
            I => \pc_rx.r_Bit_Index_1\
        );

    \I__2782\ : CEMux
    port map (
            O => \N__13900\,
            I => \N__13897\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__13897\,
            I => n5482
        );

    \I__2780\ : SRMux
    port map (
            O => \N__13894\,
            I => \N__13891\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__13891\,
            I => \N__13888\
        );

    \I__2778\ : Span4Mux_v
    port map (
            O => \N__13888\,
            I => \N__13885\
        );

    \I__2777\ : Span4Mux_h
    port map (
            O => \N__13885\,
            I => \N__13882\
        );

    \I__2776\ : Odrv4
    port map (
            O => \N__13882\,
            I => \pc_rx.n2676\
        );

    \I__2775\ : InMux
    port map (
            O => \N__13879\,
            I => \N__13874\
        );

    \I__2774\ : InMux
    port map (
            O => \N__13878\,
            I => \N__13869\
        );

    \I__2773\ : InMux
    port map (
            O => \N__13877\,
            I => \N__13869\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__13874\,
            I => debug_led3
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__13869\,
            I => debug_led3
        );

    \I__2770\ : InMux
    port map (
            O => \N__13864\,
            I => \N__13861\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__13861\,
            I => uart_rx_complete_prev
        );

    \I__2768\ : InMux
    port map (
            O => \N__13858\,
            I => \N__13855\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__13855\,
            I => \bluejay_data_inst.n19\
        );

    \I__2766\ : InMux
    port map (
            O => \N__13852\,
            I => \N__13849\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__13849\,
            I => \N__13845\
        );

    \I__2764\ : InMux
    port map (
            O => \N__13848\,
            I => \N__13842\
        );

    \I__2763\ : Odrv4
    port map (
            O => \N__13845\,
            I => n4_adj_666
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__13842\,
            I => n4_adj_666
        );

    \I__2761\ : InMux
    port map (
            O => \N__13837\,
            I => \N__13834\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__13834\,
            I => \N__13829\
        );

    \I__2759\ : InMux
    port map (
            O => \N__13833\,
            I => \N__13826\
        );

    \I__2758\ : InMux
    port map (
            O => \N__13832\,
            I => \N__13823\
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__13829\,
            I => n2471
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__13826\,
            I => n2471
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__13823\,
            I => n2471
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__13816\,
            I => \N__13812\
        );

    \I__2753\ : InMux
    port map (
            O => \N__13815\,
            I => \N__13807\
        );

    \I__2752\ : InMux
    port map (
            O => \N__13812\,
            I => \N__13807\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__13807\,
            I => pc_data_rx_2
        );

    \I__2750\ : CascadeMux
    port map (
            O => \N__13804\,
            I => \N__13801\
        );

    \I__2749\ : InMux
    port map (
            O => \N__13801\,
            I => \N__13797\
        );

    \I__2748\ : InMux
    port map (
            O => \N__13800\,
            I => \N__13794\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__13797\,
            I => \N__13788\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__13794\,
            I => \N__13788\
        );

    \I__2745\ : InMux
    port map (
            O => \N__13793\,
            I => \N__13785\
        );

    \I__2744\ : Span4Mux_h
    port map (
            O => \N__13788\,
            I => \N__13782\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__13785\,
            I => tx_data_byte_2
        );

    \I__2742\ : Odrv4
    port map (
            O => \N__13782\,
            I => tx_data_byte_2
        );

    \I__2741\ : CascadeMux
    port map (
            O => \N__13777\,
            I => \N__13774\
        );

    \I__2740\ : InMux
    port map (
            O => \N__13774\,
            I => \N__13771\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__13771\,
            I => \N__13767\
        );

    \I__2738\ : InMux
    port map (
            O => \N__13770\,
            I => \N__13764\
        );

    \I__2737\ : Span4Mux_v
    port map (
            O => \N__13767\,
            I => \N__13760\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__13764\,
            I => \N__13757\
        );

    \I__2735\ : InMux
    port map (
            O => \N__13763\,
            I => \N__13754\
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__13760\,
            I => tx_data_byte_3
        );

    \I__2733\ : Odrv4
    port map (
            O => \N__13757\,
            I => tx_data_byte_3
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__13754\,
            I => tx_data_byte_3
        );

    \I__2731\ : InMux
    port map (
            O => \N__13747\,
            I => \N__13744\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__13744\,
            I => \N__13741\
        );

    \I__2729\ : Span4Mux_v
    port map (
            O => \N__13741\,
            I => \N__13737\
        );

    \I__2728\ : InMux
    port map (
            O => \N__13740\,
            I => \N__13734\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__13737\,
            I => tx_addr_byte_3
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__13734\,
            I => tx_addr_byte_3
        );

    \I__2725\ : InMux
    port map (
            O => \N__13729\,
            I => \N__13726\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__13726\,
            I => \N__13723\
        );

    \I__2723\ : Span4Mux_v
    port map (
            O => \N__13723\,
            I => \N__13718\
        );

    \I__2722\ : InMux
    port map (
            O => \N__13722\,
            I => \N__13715\
        );

    \I__2721\ : InMux
    port map (
            O => \N__13721\,
            I => \N__13712\
        );

    \I__2720\ : Odrv4
    port map (
            O => \N__13718\,
            I => tx_data_byte_0
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__13715\,
            I => tx_data_byte_0
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__13712\,
            I => tx_data_byte_0
        );

    \I__2717\ : InMux
    port map (
            O => \N__13705\,
            I => \N__13702\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__13702\,
            I => \N__13699\
        );

    \I__2715\ : Span4Mux_v
    port map (
            O => \N__13699\,
            I => \N__13695\
        );

    \I__2714\ : InMux
    port map (
            O => \N__13698\,
            I => \N__13692\
        );

    \I__2713\ : Odrv4
    port map (
            O => \N__13695\,
            I => tx_addr_byte_0
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__13692\,
            I => tx_addr_byte_0
        );

    \I__2711\ : InMux
    port map (
            O => \N__13687\,
            I => \N__13684\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__13684\,
            I => \bluejay_data_inst.n5531\
        );

    \I__2709\ : InMux
    port map (
            O => \N__13681\,
            I => \N__13676\
        );

    \I__2708\ : InMux
    port map (
            O => \N__13680\,
            I => \N__13673\
        );

    \I__2707\ : InMux
    port map (
            O => \N__13679\,
            I => \N__13670\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__13676\,
            I => \pc_rx.r_Clock_Count_1\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__13673\,
            I => \pc_rx.r_Clock_Count_1\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__13670\,
            I => \pc_rx.r_Clock_Count_1\
        );

    \I__2703\ : InMux
    port map (
            O => \N__13663\,
            I => \N__13658\
        );

    \I__2702\ : InMux
    port map (
            O => \N__13662\,
            I => \N__13655\
        );

    \I__2701\ : InMux
    port map (
            O => \N__13661\,
            I => \N__13652\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__13658\,
            I => \pc_rx.r_Clock_Count_4\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__13655\,
            I => \pc_rx.r_Clock_Count_4\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__13652\,
            I => \pc_rx.r_Clock_Count_4\
        );

    \I__2697\ : InMux
    port map (
            O => \N__13645\,
            I => \N__13640\
        );

    \I__2696\ : InMux
    port map (
            O => \N__13644\,
            I => \N__13637\
        );

    \I__2695\ : InMux
    port map (
            O => \N__13643\,
            I => \N__13634\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__13640\,
            I => \pc_rx.r_Clock_Count_0\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__13637\,
            I => \pc_rx.r_Clock_Count_0\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__13634\,
            I => \pc_rx.r_Clock_Count_0\
        );

    \I__2691\ : InMux
    port map (
            O => \N__13627\,
            I => \N__13624\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__13624\,
            I => \pc_rx.n4\
        );

    \I__2689\ : InMux
    port map (
            O => \N__13621\,
            I => \N__13618\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__13618\,
            I => \N__13614\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__13617\,
            I => \N__13611\
        );

    \I__2686\ : Span4Mux_h
    port map (
            O => \N__13614\,
            I => \N__13608\
        );

    \I__2685\ : InMux
    port map (
            O => \N__13611\,
            I => \N__13605\
        );

    \I__2684\ : Odrv4
    port map (
            O => \N__13608\,
            I => pc_data_rx_0
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__13605\,
            I => pc_data_rx_0
        );

    \I__2682\ : CascadeMux
    port map (
            O => \N__13600\,
            I => \usb_to_bluejay_if_inst.n5438_cascade_\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__13597\,
            I => \N__13594\
        );

    \I__2680\ : InMux
    port map (
            O => \N__13594\,
            I => \N__13591\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__13591\,
            I => \N__13588\
        );

    \I__2678\ : Span4Mux_h
    port map (
            O => \N__13588\,
            I => \N__13585\
        );

    \I__2677\ : Span4Mux_v
    port map (
            O => \N__13585\,
            I => \N__13581\
        );

    \I__2676\ : InMux
    port map (
            O => \N__13584\,
            I => \N__13578\
        );

    \I__2675\ : Odrv4
    port map (
            O => \N__13581\,
            I => tx_addr_byte_6
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__13578\,
            I => tx_addr_byte_6
        );

    \I__2673\ : InMux
    port map (
            O => \N__13573\,
            I => \N__13570\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__13570\,
            I => \N__13566\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__13569\,
            I => \N__13563\
        );

    \I__2670\ : Span4Mux_h
    port map (
            O => \N__13566\,
            I => \N__13559\
        );

    \I__2669\ : InMux
    port map (
            O => \N__13563\,
            I => \N__13554\
        );

    \I__2668\ : InMux
    port map (
            O => \N__13562\,
            I => \N__13554\
        );

    \I__2667\ : Odrv4
    port map (
            O => \N__13559\,
            I => tx_data_byte_6
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__13554\,
            I => tx_data_byte_6
        );

    \I__2665\ : InMux
    port map (
            O => \N__13549\,
            I => \N__13545\
        );

    \I__2664\ : InMux
    port map (
            O => \N__13548\,
            I => \N__13542\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__13545\,
            I => \N__13539\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__13542\,
            I => n3672
        );

    \I__2661\ : Odrv4
    port map (
            O => \N__13539\,
            I => n3672
        );

    \I__2660\ : CascadeMux
    port map (
            O => \N__13534\,
            I => \N__13530\
        );

    \I__2659\ : InMux
    port map (
            O => \N__13533\,
            I => \N__13525\
        );

    \I__2658\ : InMux
    port map (
            O => \N__13530\,
            I => \N__13525\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__13525\,
            I => pc_data_rx_6
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__13522\,
            I => \pc_rx.n5522_cascade_\
        );

    \I__2655\ : CascadeMux
    port map (
            O => \N__13519\,
            I => \n5482_cascade_\
        );

    \I__2654\ : InMux
    port map (
            O => \N__13516\,
            I => \N__13511\
        );

    \I__2653\ : InMux
    port map (
            O => \N__13515\,
            I => \N__13506\
        );

    \I__2652\ : InMux
    port map (
            O => \N__13514\,
            I => \N__13506\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__13511\,
            I => n3753
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__13506\,
            I => n3753
        );

    \I__2649\ : InMux
    port map (
            O => \N__13501\,
            I => \N__13498\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__13498\,
            I => \N__13489\
        );

    \I__2647\ : InMux
    port map (
            O => \N__13497\,
            I => \N__13486\
        );

    \I__2646\ : InMux
    port map (
            O => \N__13496\,
            I => \N__13481\
        );

    \I__2645\ : InMux
    port map (
            O => \N__13495\,
            I => \N__13481\
        );

    \I__2644\ : InMux
    port map (
            O => \N__13494\,
            I => \N__13474\
        );

    \I__2643\ : InMux
    port map (
            O => \N__13493\,
            I => \N__13474\
        );

    \I__2642\ : InMux
    port map (
            O => \N__13492\,
            I => \N__13474\
        );

    \I__2641\ : Odrv4
    port map (
            O => \N__13489\,
            I => \r_SM_Main_2_N_246_2\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__13486\,
            I => \r_SM_Main_2_N_246_2\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__13481\,
            I => \r_SM_Main_2_N_246_2\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__13474\,
            I => \r_SM_Main_2_N_246_2\
        );

    \I__2637\ : InMux
    port map (
            O => \N__13465\,
            I => \N__13450\
        );

    \I__2636\ : InMux
    port map (
            O => \N__13464\,
            I => \N__13450\
        );

    \I__2635\ : InMux
    port map (
            O => \N__13463\,
            I => \N__13450\
        );

    \I__2634\ : InMux
    port map (
            O => \N__13462\,
            I => \N__13450\
        );

    \I__2633\ : InMux
    port map (
            O => \N__13461\,
            I => \N__13443\
        );

    \I__2632\ : InMux
    port map (
            O => \N__13460\,
            I => \N__13438\
        );

    \I__2631\ : InMux
    port map (
            O => \N__13459\,
            I => \N__13438\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__13450\,
            I => \N__13435\
        );

    \I__2629\ : InMux
    port map (
            O => \N__13449\,
            I => \N__13432\
        );

    \I__2628\ : InMux
    port map (
            O => \N__13448\,
            I => \N__13427\
        );

    \I__2627\ : InMux
    port map (
            O => \N__13447\,
            I => \N__13427\
        );

    \I__2626\ : InMux
    port map (
            O => \N__13446\,
            I => \N__13424\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__13443\,
            I => \N__13421\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__13438\,
            I => \N__13418\
        );

    \I__2623\ : Span4Mux_h
    port map (
            O => \N__13435\,
            I => \N__13415\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__13432\,
            I => \r_SM_Main_0\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__13427\,
            I => \r_SM_Main_0\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__13424\,
            I => \r_SM_Main_0\
        );

    \I__2619\ : Odrv4
    port map (
            O => \N__13421\,
            I => \r_SM_Main_0\
        );

    \I__2618\ : Odrv12
    port map (
            O => \N__13418\,
            I => \r_SM_Main_0\
        );

    \I__2617\ : Odrv4
    port map (
            O => \N__13415\,
            I => \r_SM_Main_0\
        );

    \I__2616\ : InMux
    port map (
            O => \N__13402\,
            I => \N__13394\
        );

    \I__2615\ : InMux
    port map (
            O => \N__13401\,
            I => \N__13394\
        );

    \I__2614\ : SRMux
    port map (
            O => \N__13400\,
            I => \N__13386\
        );

    \I__2613\ : InMux
    port map (
            O => \N__13399\,
            I => \N__13383\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__13394\,
            I => \N__13380\
        );

    \I__2611\ : InMux
    port map (
            O => \N__13393\,
            I => \N__13371\
        );

    \I__2610\ : InMux
    port map (
            O => \N__13392\,
            I => \N__13371\
        );

    \I__2609\ : InMux
    port map (
            O => \N__13391\,
            I => \N__13371\
        );

    \I__2608\ : InMux
    port map (
            O => \N__13390\,
            I => \N__13371\
        );

    \I__2607\ : InMux
    port map (
            O => \N__13389\,
            I => \N__13368\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__13386\,
            I => \r_SM_Main_2\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__13383\,
            I => \r_SM_Main_2\
        );

    \I__2604\ : Odrv4
    port map (
            O => \N__13380\,
            I => \r_SM_Main_2\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__13371\,
            I => \r_SM_Main_2\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__13368\,
            I => \r_SM_Main_2\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__13357\,
            I => \n2502_cascade_\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__13354\,
            I => \N__13349\
        );

    \I__2599\ : CascadeMux
    port map (
            O => \N__13353\,
            I => \N__13344\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__13352\,
            I => \N__13341\
        );

    \I__2597\ : InMux
    port map (
            O => \N__13349\,
            I => \N__13333\
        );

    \I__2596\ : InMux
    port map (
            O => \N__13348\,
            I => \N__13330\
        );

    \I__2595\ : InMux
    port map (
            O => \N__13347\,
            I => \N__13321\
        );

    \I__2594\ : InMux
    port map (
            O => \N__13344\,
            I => \N__13321\
        );

    \I__2593\ : InMux
    port map (
            O => \N__13341\,
            I => \N__13321\
        );

    \I__2592\ : InMux
    port map (
            O => \N__13340\,
            I => \N__13321\
        );

    \I__2591\ : CascadeMux
    port map (
            O => \N__13339\,
            I => \N__13318\
        );

    \I__2590\ : InMux
    port map (
            O => \N__13338\,
            I => \N__13312\
        );

    \I__2589\ : InMux
    port map (
            O => \N__13337\,
            I => \N__13312\
        );

    \I__2588\ : InMux
    port map (
            O => \N__13336\,
            I => \N__13309\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__13333\,
            I => \N__13302\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__13330\,
            I => \N__13302\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__13321\,
            I => \N__13302\
        );

    \I__2584\ : InMux
    port map (
            O => \N__13318\,
            I => \N__13299\
        );

    \I__2583\ : InMux
    port map (
            O => \N__13317\,
            I => \N__13296\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__13312\,
            I => \N__13293\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__13309\,
            I => \N__13290\
        );

    \I__2580\ : Span4Mux_h
    port map (
            O => \N__13302\,
            I => \N__13287\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__13299\,
            I => \r_SM_Main_1\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__13296\,
            I => \r_SM_Main_1\
        );

    \I__2577\ : Odrv12
    port map (
            O => \N__13293\,
            I => \r_SM_Main_1\
        );

    \I__2576\ : Odrv4
    port map (
            O => \N__13290\,
            I => \r_SM_Main_1\
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__13287\,
            I => \r_SM_Main_1\
        );

    \I__2574\ : CascadeMux
    port map (
            O => \N__13276\,
            I => \bluejay_data_inst.n1041_cascade_\
        );

    \I__2573\ : CascadeMux
    port map (
            O => \N__13273\,
            I => \bluejay_data_inst.state_timeout_counter_7_N_122_2_cascade_\
        );

    \I__2572\ : CascadeMux
    port map (
            O => \N__13270\,
            I => \bluejay_data_inst.n18_cascade_\
        );

    \I__2571\ : InMux
    port map (
            O => \N__13267\,
            I => \N__13264\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__13264\,
            I => \bluejay_data_inst.n20\
        );

    \I__2569\ : InMux
    port map (
            O => \N__13261\,
            I => \N__13256\
        );

    \I__2568\ : InMux
    port map (
            O => \N__13260\,
            I => \N__13251\
        );

    \I__2567\ : InMux
    port map (
            O => \N__13259\,
            I => \N__13251\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__13256\,
            I => \bluejay_data_inst.n1675\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__13251\,
            I => \bluejay_data_inst.n1675\
        );

    \I__2564\ : InMux
    port map (
            O => \N__13246\,
            I => \N__13243\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__13243\,
            I => \N__13240\
        );

    \I__2562\ : Span12Mux_h
    port map (
            O => \N__13240\,
            I => \N__13237\
        );

    \I__2561\ : Span12Mux_v
    port map (
            O => \N__13237\,
            I => \N__13234\
        );

    \I__2560\ : Odrv12
    port map (
            O => \N__13234\,
            I => \FIFO_D1_c_1\
        );

    \I__2559\ : IoInMux
    port map (
            O => \N__13231\,
            I => \N__13228\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__13228\,
            I => \N__13225\
        );

    \I__2557\ : Span4Mux_s3_v
    port map (
            O => \N__13225\,
            I => \N__13222\
        );

    \I__2556\ : Sp12to4
    port map (
            O => \N__13222\,
            I => \N__13219\
        );

    \I__2555\ : Span12Mux_s10_h
    port map (
            O => \N__13219\,
            I => \N__13216\
        );

    \I__2554\ : Span12Mux_v
    port map (
            O => \N__13216\,
            I => \N__13213\
        );

    \I__2553\ : Odrv12
    port map (
            O => \N__13213\,
            I => \DATA1_c_1\
        );

    \I__2552\ : InMux
    port map (
            O => \N__13210\,
            I => \N__13207\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__13207\,
            I => \N__13204\
        );

    \I__2550\ : Span4Mux_v
    port map (
            O => \N__13204\,
            I => \N__13201\
        );

    \I__2549\ : Sp12to4
    port map (
            O => \N__13201\,
            I => \N__13198\
        );

    \I__2548\ : Span12Mux_h
    port map (
            O => \N__13198\,
            I => \N__13195\
        );

    \I__2547\ : Span12Mux_v
    port map (
            O => \N__13195\,
            I => \N__13192\
        );

    \I__2546\ : Odrv12
    port map (
            O => \N__13192\,
            I => \FIFO_D21_c_21\
        );

    \I__2545\ : IoInMux
    port map (
            O => \N__13189\,
            I => \N__13186\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__13186\,
            I => \N__13183\
        );

    \I__2543\ : IoSpan4Mux
    port map (
            O => \N__13183\,
            I => \N__13180\
        );

    \I__2542\ : Span4Mux_s2_v
    port map (
            O => \N__13180\,
            I => \N__13177\
        );

    \I__2541\ : Sp12to4
    port map (
            O => \N__13177\,
            I => \N__13174\
        );

    \I__2540\ : Span12Mux_h
    port map (
            O => \N__13174\,
            I => \N__13171\
        );

    \I__2539\ : Odrv12
    port map (
            O => \N__13171\,
            I => \DATA21_c_21\
        );

    \I__2538\ : InMux
    port map (
            O => \N__13168\,
            I => \N__13163\
        );

    \I__2537\ : InMux
    port map (
            O => \N__13167\,
            I => \N__13160\
        );

    \I__2536\ : InMux
    port map (
            O => \N__13166\,
            I => \N__13157\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__13163\,
            I => \pc_rx.r_Clock_Count_7\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__13160\,
            I => \pc_rx.r_Clock_Count_7\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__13157\,
            I => \pc_rx.r_Clock_Count_7\
        );

    \I__2532\ : InMux
    port map (
            O => \N__13150\,
            I => \pc_rx.n4813\
        );

    \I__2531\ : InMux
    port map (
            O => \N__13147\,
            I => \N__13143\
        );

    \I__2530\ : InMux
    port map (
            O => \N__13146\,
            I => \N__13139\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__13143\,
            I => \N__13136\
        );

    \I__2528\ : InMux
    port map (
            O => \N__13142\,
            I => \N__13133\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__13139\,
            I => \pc_rx.r_Clock_Count_8\
        );

    \I__2526\ : Odrv4
    port map (
            O => \N__13136\,
            I => \pc_rx.r_Clock_Count_8\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__13133\,
            I => \pc_rx.r_Clock_Count_8\
        );

    \I__2524\ : InMux
    port map (
            O => \N__13126\,
            I => \bfn_13_7_0_\
        );

    \I__2523\ : InMux
    port map (
            O => \N__13123\,
            I => \pc_rx.n4815\
        );

    \I__2522\ : InMux
    port map (
            O => \N__13120\,
            I => \N__13115\
        );

    \I__2521\ : InMux
    port map (
            O => \N__13119\,
            I => \N__13112\
        );

    \I__2520\ : InMux
    port map (
            O => \N__13118\,
            I => \N__13109\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__13115\,
            I => \N__13106\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__13112\,
            I => \pc_rx.r_Clock_Count_9\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__13109\,
            I => \pc_rx.r_Clock_Count_9\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__13106\,
            I => \pc_rx.r_Clock_Count_9\
        );

    \I__2515\ : CEMux
    port map (
            O => \N__13099\,
            I => \N__13096\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__13096\,
            I => \N__13092\
        );

    \I__2513\ : CEMux
    port map (
            O => \N__13095\,
            I => \N__13089\
        );

    \I__2512\ : Span4Mux_h
    port map (
            O => \N__13092\,
            I => \N__13086\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__13089\,
            I => \N__13083\
        );

    \I__2510\ : Odrv4
    port map (
            O => \N__13086\,
            I => \pc_rx.n2566\
        );

    \I__2509\ : Odrv4
    port map (
            O => \N__13083\,
            I => \pc_rx.n2566\
        );

    \I__2508\ : SRMux
    port map (
            O => \N__13078\,
            I => \N__13074\
        );

    \I__2507\ : SRMux
    port map (
            O => \N__13077\,
            I => \N__13071\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__13074\,
            I => \N__13068\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__13071\,
            I => \N__13065\
        );

    \I__2504\ : Span4Mux_h
    port map (
            O => \N__13068\,
            I => \N__13062\
        );

    \I__2503\ : Span4Mux_h
    port map (
            O => \N__13065\,
            I => \N__13059\
        );

    \I__2502\ : Odrv4
    port map (
            O => \N__13062\,
            I => \pc_rx.n2705\
        );

    \I__2501\ : Odrv4
    port map (
            O => \N__13059\,
            I => \pc_rx.n2705\
        );

    \I__2500\ : InMux
    port map (
            O => \N__13054\,
            I => \N__13047\
        );

    \I__2499\ : InMux
    port map (
            O => \N__13053\,
            I => \N__13044\
        );

    \I__2498\ : InMux
    port map (
            O => \N__13052\,
            I => \N__13040\
        );

    \I__2497\ : InMux
    port map (
            O => \N__13051\,
            I => \N__13025\
        );

    \I__2496\ : InMux
    port map (
            O => \N__13050\,
            I => \N__13025\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__13047\,
            I => \N__13022\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__13044\,
            I => \N__13019\
        );

    \I__2493\ : InMux
    port map (
            O => \N__13043\,
            I => \N__13016\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__13040\,
            I => \N__13013\
        );

    \I__2491\ : InMux
    port map (
            O => \N__13039\,
            I => \N__13004\
        );

    \I__2490\ : InMux
    port map (
            O => \N__13038\,
            I => \N__13004\
        );

    \I__2489\ : InMux
    port map (
            O => \N__13037\,
            I => \N__13004\
        );

    \I__2488\ : InMux
    port map (
            O => \N__13036\,
            I => \N__13004\
        );

    \I__2487\ : InMux
    port map (
            O => \N__13035\,
            I => \N__13001\
        );

    \I__2486\ : InMux
    port map (
            O => \N__13034\,
            I => \N__12998\
        );

    \I__2485\ : InMux
    port map (
            O => \N__13033\,
            I => \N__12989\
        );

    \I__2484\ : InMux
    port map (
            O => \N__13032\,
            I => \N__12989\
        );

    \I__2483\ : InMux
    port map (
            O => \N__13031\,
            I => \N__12989\
        );

    \I__2482\ : InMux
    port map (
            O => \N__13030\,
            I => \N__12989\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__13025\,
            I => state_reg_2
        );

    \I__2480\ : Odrv12
    port map (
            O => \N__13022\,
            I => state_reg_2
        );

    \I__2479\ : Odrv4
    port map (
            O => \N__13019\,
            I => state_reg_2
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__13016\,
            I => state_reg_2
        );

    \I__2477\ : Odrv12
    port map (
            O => \N__13013\,
            I => state_reg_2
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__13004\,
            I => state_reg_2
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__13001\,
            I => state_reg_2
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__12998\,
            I => state_reg_2
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__12989\,
            I => state_reg_2
        );

    \I__2472\ : SRMux
    port map (
            O => \N__12970\,
            I => \N__12965\
        );

    \I__2471\ : InMux
    port map (
            O => \N__12969\,
            I => \N__12962\
        );

    \I__2470\ : InMux
    port map (
            O => \N__12968\,
            I => \N__12957\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__12965\,
            I => \N__12954\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__12962\,
            I => \N__12951\
        );

    \I__2467\ : InMux
    port map (
            O => \N__12961\,
            I => \N__12946\
        );

    \I__2466\ : InMux
    port map (
            O => \N__12960\,
            I => \N__12946\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__12957\,
            I => \N__12934\
        );

    \I__2464\ : Span4Mux_h
    port map (
            O => \N__12954\,
            I => \N__12914\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__12951\,
            I => \N__12911\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__12946\,
            I => \N__12908\
        );

    \I__2461\ : InMux
    port map (
            O => \N__12945\,
            I => \N__12905\
        );

    \I__2460\ : InMux
    port map (
            O => \N__12944\,
            I => \N__12888\
        );

    \I__2459\ : InMux
    port map (
            O => \N__12943\,
            I => \N__12888\
        );

    \I__2458\ : InMux
    port map (
            O => \N__12942\,
            I => \N__12888\
        );

    \I__2457\ : InMux
    port map (
            O => \N__12941\,
            I => \N__12888\
        );

    \I__2456\ : InMux
    port map (
            O => \N__12940\,
            I => \N__12888\
        );

    \I__2455\ : InMux
    port map (
            O => \N__12939\,
            I => \N__12888\
        );

    \I__2454\ : InMux
    port map (
            O => \N__12938\,
            I => \N__12888\
        );

    \I__2453\ : InMux
    port map (
            O => \N__12937\,
            I => \N__12888\
        );

    \I__2452\ : Span4Mux_v
    port map (
            O => \N__12934\,
            I => \N__12885\
        );

    \I__2451\ : InMux
    port map (
            O => \N__12933\,
            I => \N__12874\
        );

    \I__2450\ : InMux
    port map (
            O => \N__12932\,
            I => \N__12874\
        );

    \I__2449\ : InMux
    port map (
            O => \N__12931\,
            I => \N__12874\
        );

    \I__2448\ : InMux
    port map (
            O => \N__12930\,
            I => \N__12874\
        );

    \I__2447\ : InMux
    port map (
            O => \N__12929\,
            I => \N__12874\
        );

    \I__2446\ : InMux
    port map (
            O => \N__12928\,
            I => \N__12865\
        );

    \I__2445\ : InMux
    port map (
            O => \N__12927\,
            I => \N__12865\
        );

    \I__2444\ : InMux
    port map (
            O => \N__12926\,
            I => \N__12865\
        );

    \I__2443\ : InMux
    port map (
            O => \N__12925\,
            I => \N__12865\
        );

    \I__2442\ : InMux
    port map (
            O => \N__12924\,
            I => \N__12862\
        );

    \I__2441\ : InMux
    port map (
            O => \N__12923\,
            I => \N__12859\
        );

    \I__2440\ : InMux
    port map (
            O => \N__12922\,
            I => \N__12846\
        );

    \I__2439\ : InMux
    port map (
            O => \N__12921\,
            I => \N__12846\
        );

    \I__2438\ : InMux
    port map (
            O => \N__12920\,
            I => \N__12846\
        );

    \I__2437\ : InMux
    port map (
            O => \N__12919\,
            I => \N__12846\
        );

    \I__2436\ : InMux
    port map (
            O => \N__12918\,
            I => \N__12846\
        );

    \I__2435\ : InMux
    port map (
            O => \N__12917\,
            I => \N__12846\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__12914\,
            I => state_reg_1
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__12911\,
            I => state_reg_1
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__12908\,
            I => state_reg_1
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__12905\,
            I => state_reg_1
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__12888\,
            I => state_reg_1
        );

    \I__2429\ : Odrv4
    port map (
            O => \N__12885\,
            I => state_reg_1
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__12874\,
            I => state_reg_1
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__12865\,
            I => state_reg_1
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__12862\,
            I => state_reg_1
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__12859\,
            I => state_reg_1
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__12846\,
            I => state_reg_1
        );

    \I__2423\ : InMux
    port map (
            O => \N__12823\,
            I => \N__12820\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__12820\,
            I => \N__12817\
        );

    \I__2421\ : Span4Mux_h
    port map (
            O => \N__12817\,
            I => \N__12814\
        );

    \I__2420\ : Odrv4
    port map (
            O => \N__12814\,
            I => tx_shift_reg_0
        );

    \I__2419\ : SRMux
    port map (
            O => \N__12811\,
            I => \N__12808\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__12808\,
            I => \N__12805\
        );

    \I__2417\ : Span4Mux_h
    port map (
            O => \N__12805\,
            I => \N__12802\
        );

    \I__2416\ : Span4Mux_h
    port map (
            O => \N__12802\,
            I => \N__12799\
        );

    \I__2415\ : Odrv4
    port map (
            O => \N__12799\,
            I => n989
        );

    \I__2414\ : CascadeMux
    port map (
            O => \N__12796\,
            I => \bluejay_data_inst.n1040_cascade_\
        );

    \I__2413\ : CascadeMux
    port map (
            O => \N__12793\,
            I => \bluejay_data_inst.state_timeout_counter_7_N_122_3_cascade_\
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__12790\,
            I => \bluejay_data_inst.n8_adj_656_cascade_\
        );

    \I__2411\ : InMux
    port map (
            O => \N__12787\,
            I => \N__12784\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__12784\,
            I => \bluejay_data_inst.state_timeout_counter_7_N_122_3\
        );

    \I__2409\ : CascadeMux
    port map (
            O => \N__12781\,
            I => \pc_rx.n2429_cascade_\
        );

    \I__2408\ : InMux
    port map (
            O => \N__12778\,
            I => \bfn_13_6_0_\
        );

    \I__2407\ : InMux
    port map (
            O => \N__12775\,
            I => \pc_rx.n4807\
        );

    \I__2406\ : InMux
    port map (
            O => \N__12772\,
            I => \N__12767\
        );

    \I__2405\ : InMux
    port map (
            O => \N__12771\,
            I => \N__12764\
        );

    \I__2404\ : InMux
    port map (
            O => \N__12770\,
            I => \N__12761\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__12767\,
            I => \pc_rx.r_Clock_Count_2\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__12764\,
            I => \pc_rx.r_Clock_Count_2\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__12761\,
            I => \pc_rx.r_Clock_Count_2\
        );

    \I__2400\ : InMux
    port map (
            O => \N__12754\,
            I => \pc_rx.n4808\
        );

    \I__2399\ : InMux
    port map (
            O => \N__12751\,
            I => \N__12746\
        );

    \I__2398\ : InMux
    port map (
            O => \N__12750\,
            I => \N__12743\
        );

    \I__2397\ : InMux
    port map (
            O => \N__12749\,
            I => \N__12740\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__12746\,
            I => \pc_rx.r_Clock_Count_3\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__12743\,
            I => \pc_rx.r_Clock_Count_3\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__12740\,
            I => \pc_rx.r_Clock_Count_3\
        );

    \I__2393\ : InMux
    port map (
            O => \N__12733\,
            I => \pc_rx.n4809\
        );

    \I__2392\ : InMux
    port map (
            O => \N__12730\,
            I => \pc_rx.n4810\
        );

    \I__2391\ : InMux
    port map (
            O => \N__12727\,
            I => \N__12722\
        );

    \I__2390\ : InMux
    port map (
            O => \N__12726\,
            I => \N__12719\
        );

    \I__2389\ : InMux
    port map (
            O => \N__12725\,
            I => \N__12716\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__12722\,
            I => \pc_rx.r_Clock_Count_5\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__12719\,
            I => \pc_rx.r_Clock_Count_5\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__12716\,
            I => \pc_rx.r_Clock_Count_5\
        );

    \I__2385\ : InMux
    port map (
            O => \N__12709\,
            I => \pc_rx.n4811\
        );

    \I__2384\ : InMux
    port map (
            O => \N__12706\,
            I => \N__12701\
        );

    \I__2383\ : InMux
    port map (
            O => \N__12705\,
            I => \N__12698\
        );

    \I__2382\ : InMux
    port map (
            O => \N__12704\,
            I => \N__12695\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__12701\,
            I => \pc_rx.r_Clock_Count_6\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__12698\,
            I => \pc_rx.r_Clock_Count_6\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__12695\,
            I => \pc_rx.r_Clock_Count_6\
        );

    \I__2378\ : InMux
    port map (
            O => \N__12688\,
            I => \pc_rx.n4812\
        );

    \I__2377\ : InMux
    port map (
            O => \N__12685\,
            I => \N__12682\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__12682\,
            I => n2468
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__12679\,
            I => \N__12675\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__12678\,
            I => \N__12672\
        );

    \I__2373\ : InMux
    port map (
            O => \N__12675\,
            I => \N__12667\
        );

    \I__2372\ : InMux
    port map (
            O => \N__12672\,
            I => \N__12667\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__12667\,
            I => pc_data_rx_4
        );

    \I__2370\ : InMux
    port map (
            O => \N__12664\,
            I => \N__12661\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__12661\,
            I => \pc_rx.n3803\
        );

    \I__2368\ : CascadeMux
    port map (
            O => \N__12658\,
            I => \n2475_cascade_\
        );

    \I__2367\ : InMux
    port map (
            O => \N__12655\,
            I => \N__12651\
        );

    \I__2366\ : InMux
    port map (
            O => \N__12654\,
            I => \N__12648\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__12651\,
            I => pc_data_rx_7
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__12648\,
            I => pc_data_rx_7
        );

    \I__2363\ : InMux
    port map (
            O => \N__12643\,
            I => \N__12639\
        );

    \I__2362\ : InMux
    port map (
            O => \N__12642\,
            I => \N__12636\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__12639\,
            I => n2475
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__12636\,
            I => n2475
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__12631\,
            I => \N__12627\
        );

    \I__2358\ : InMux
    port map (
            O => \N__12630\,
            I => \N__12624\
        );

    \I__2357\ : InMux
    port map (
            O => \N__12627\,
            I => \N__12621\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__12624\,
            I => pc_data_rx_3
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__12621\,
            I => pc_data_rx_3
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__12616\,
            I => \pc_rx.n2465_cascade_\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__12613\,
            I => \pc_rx.n4887_cascade_\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__12610\,
            I => \r_SM_Main_2_N_246_2_cascade_\
        );

    \I__2351\ : InMux
    port map (
            O => \N__12607\,
            I => \N__12603\
        );

    \I__2350\ : InMux
    port map (
            O => \N__12606\,
            I => \N__12600\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__12603\,
            I => \pc_rx.n2429\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__12600\,
            I => \pc_rx.n2429\
        );

    \I__2347\ : InMux
    port map (
            O => \N__12595\,
            I => \N__12592\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__12592\,
            I => \N__12589\
        );

    \I__2345\ : Span12Mux_v
    port map (
            O => \N__12589\,
            I => \N__12586\
        );

    \I__2344\ : Span12Mux_h
    port map (
            O => \N__12586\,
            I => \N__12583\
        );

    \I__2343\ : Odrv12
    port map (
            O => \N__12583\,
            I => \FIFO_D24_c_24\
        );

    \I__2342\ : IoInMux
    port map (
            O => \N__12580\,
            I => \N__12577\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__12577\,
            I => \N__12574\
        );

    \I__2340\ : Span4Mux_s3_v
    port map (
            O => \N__12574\,
            I => \N__12571\
        );

    \I__2339\ : Sp12to4
    port map (
            O => \N__12571\,
            I => \N__12568\
        );

    \I__2338\ : Span12Mux_h
    port map (
            O => \N__12568\,
            I => \N__12565\
        );

    \I__2337\ : Span12Mux_v
    port map (
            O => \N__12565\,
            I => \N__12562\
        );

    \I__2336\ : Odrv12
    port map (
            O => \N__12562\,
            I => \DATA24_c_24\
        );

    \I__2335\ : InMux
    port map (
            O => \N__12559\,
            I => \N__12556\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__12556\,
            I => \N__12553\
        );

    \I__2333\ : Span12Mux_v
    port map (
            O => \N__12553\,
            I => \N__12550\
        );

    \I__2332\ : Odrv12
    port map (
            O => \N__12550\,
            I => \FIFO_D5_c_5\
        );

    \I__2331\ : IoInMux
    port map (
            O => \N__12547\,
            I => \N__12544\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__12544\,
            I => \N__12541\
        );

    \I__2329\ : Span4Mux_s2_v
    port map (
            O => \N__12541\,
            I => \N__12538\
        );

    \I__2328\ : Sp12to4
    port map (
            O => \N__12538\,
            I => \N__12535\
        );

    \I__2327\ : Span12Mux_h
    port map (
            O => \N__12535\,
            I => \N__12532\
        );

    \I__2326\ : Span12Mux_v
    port map (
            O => \N__12532\,
            I => \N__12529\
        );

    \I__2325\ : Odrv12
    port map (
            O => \N__12529\,
            I => \DATA5_c_5\
        );

    \I__2324\ : InMux
    port map (
            O => \N__12526\,
            I => \N__12523\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__12523\,
            I => \N__12520\
        );

    \I__2322\ : Span12Mux_v
    port map (
            O => \N__12520\,
            I => \N__12517\
        );

    \I__2321\ : Odrv12
    port map (
            O => \N__12517\,
            I => \FIFO_D6_c_6\
        );

    \I__2320\ : IoInMux
    port map (
            O => \N__12514\,
            I => \N__12511\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__12511\,
            I => \N__12508\
        );

    \I__2318\ : IoSpan4Mux
    port map (
            O => \N__12508\,
            I => \N__12505\
        );

    \I__2317\ : Span4Mux_s3_v
    port map (
            O => \N__12505\,
            I => \N__12502\
        );

    \I__2316\ : Span4Mux_h
    port map (
            O => \N__12502\,
            I => \N__12499\
        );

    \I__2315\ : Sp12to4
    port map (
            O => \N__12499\,
            I => \N__12496\
        );

    \I__2314\ : Span12Mux_h
    port map (
            O => \N__12496\,
            I => \N__12493\
        );

    \I__2313\ : Odrv12
    port map (
            O => \N__12493\,
            I => \DATA6_c_6\
        );

    \I__2312\ : InMux
    port map (
            O => \N__12490\,
            I => \N__12484\
        );

    \I__2311\ : InMux
    port map (
            O => \N__12489\,
            I => \N__12484\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__12484\,
            I => \N__12481\
        );

    \I__2309\ : Odrv4
    port map (
            O => \N__12481\,
            I => n4
        );

    \I__2308\ : CascadeMux
    port map (
            O => \N__12478\,
            I => \N__12475\
        );

    \I__2307\ : InMux
    port map (
            O => \N__12475\,
            I => \N__12472\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__12472\,
            I => \N__12469\
        );

    \I__2305\ : Span4Mux_v
    port map (
            O => \N__12469\,
            I => \N__12464\
        );

    \I__2304\ : InMux
    port map (
            O => \N__12468\,
            I => \N__12461\
        );

    \I__2303\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12458\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__12464\,
            I => tx_data_byte_4
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__12461\,
            I => tx_data_byte_4
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__12458\,
            I => tx_data_byte_4
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__12451\,
            I => \n2468_cascade_\
        );

    \I__2298\ : InMux
    port map (
            O => \N__12448\,
            I => \N__12442\
        );

    \I__2297\ : InMux
    port map (
            O => \N__12447\,
            I => \N__12442\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__12442\,
            I => pc_data_rx_5
        );

    \I__2295\ : InMux
    port map (
            O => \N__12439\,
            I => \N__12436\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__12436\,
            I => \N__12432\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__12435\,
            I => \N__12428\
        );

    \I__2292\ : Span4Mux_v
    port map (
            O => \N__12432\,
            I => \N__12425\
        );

    \I__2291\ : InMux
    port map (
            O => \N__12431\,
            I => \N__12422\
        );

    \I__2290\ : InMux
    port map (
            O => \N__12428\,
            I => \N__12419\
        );

    \I__2289\ : Odrv4
    port map (
            O => \N__12425\,
            I => tx_data_byte_5
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__12422\,
            I => tx_data_byte_5
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__12419\,
            I => tx_data_byte_5
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__12412\,
            I => \N__12409\
        );

    \I__2285\ : InMux
    port map (
            O => \N__12409\,
            I => \N__12406\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__12406\,
            I => \tx_fifo.lscc_fifo_inst.n2\
        );

    \I__2283\ : InMux
    port map (
            O => \N__12403\,
            I => \N__12396\
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__12402\,
            I => \N__12393\
        );

    \I__2281\ : InMux
    port map (
            O => \N__12401\,
            I => \N__12386\
        );

    \I__2280\ : InMux
    port map (
            O => \N__12400\,
            I => \N__12383\
        );

    \I__2279\ : InMux
    port map (
            O => \N__12399\,
            I => \N__12374\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__12396\,
            I => \N__12371\
        );

    \I__2277\ : InMux
    port map (
            O => \N__12393\,
            I => \N__12367\
        );

    \I__2276\ : InMux
    port map (
            O => \N__12392\,
            I => \N__12358\
        );

    \I__2275\ : InMux
    port map (
            O => \N__12391\,
            I => \N__12358\
        );

    \I__2274\ : InMux
    port map (
            O => \N__12390\,
            I => \N__12358\
        );

    \I__2273\ : InMux
    port map (
            O => \N__12389\,
            I => \N__12358\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__12386\,
            I => \N__12353\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__12383\,
            I => \N__12353\
        );

    \I__2270\ : InMux
    port map (
            O => \N__12382\,
            I => \N__12350\
        );

    \I__2269\ : InMux
    port map (
            O => \N__12381\,
            I => \N__12338\
        );

    \I__2268\ : InMux
    port map (
            O => \N__12380\,
            I => \N__12338\
        );

    \I__2267\ : InMux
    port map (
            O => \N__12379\,
            I => \N__12338\
        );

    \I__2266\ : InMux
    port map (
            O => \N__12378\,
            I => \N__12338\
        );

    \I__2265\ : InMux
    port map (
            O => \N__12377\,
            I => \N__12338\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__12374\,
            I => \N__12329\
        );

    \I__2263\ : Span4Mux_h
    port map (
            O => \N__12371\,
            I => \N__12329\
        );

    \I__2262\ : InMux
    port map (
            O => \N__12370\,
            I => \N__12325\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__12367\,
            I => \N__12316\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__12358\,
            I => \N__12316\
        );

    \I__2259\ : Span4Mux_h
    port map (
            O => \N__12353\,
            I => \N__12316\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__12350\,
            I => \N__12316\
        );

    \I__2257\ : InMux
    port map (
            O => \N__12349\,
            I => \N__12313\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__12338\,
            I => \N__12310\
        );

    \I__2255\ : InMux
    port map (
            O => \N__12337\,
            I => \N__12307\
        );

    \I__2254\ : InMux
    port map (
            O => \N__12336\,
            I => \N__12302\
        );

    \I__2253\ : InMux
    port map (
            O => \N__12335\,
            I => \N__12302\
        );

    \I__2252\ : InMux
    port map (
            O => \N__12334\,
            I => \N__12299\
        );

    \I__2251\ : Span4Mux_h
    port map (
            O => \N__12329\,
            I => \N__12296\
        );

    \I__2250\ : InMux
    port map (
            O => \N__12328\,
            I => \N__12293\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__12325\,
            I => \N__12288\
        );

    \I__2248\ : Span4Mux_v
    port map (
            O => \N__12316\,
            I => \N__12288\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__12313\,
            I => rd_addr_r_1
        );

    \I__2246\ : Odrv12
    port map (
            O => \N__12310\,
            I => rd_addr_r_1
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__12307\,
            I => rd_addr_r_1
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__12302\,
            I => rd_addr_r_1
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__12299\,
            I => rd_addr_r_1
        );

    \I__2242\ : Odrv4
    port map (
            O => \N__12296\,
            I => rd_addr_r_1
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__12293\,
            I => rd_addr_r_1
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__12288\,
            I => rd_addr_r_1
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__12271\,
            I => \n32_cascade_\
        );

    \I__2238\ : InMux
    port map (
            O => \N__12268\,
            I => \N__12264\
        );

    \I__2237\ : InMux
    port map (
            O => \N__12267\,
            I => \N__12261\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__12264\,
            I => \N__12255\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__12261\,
            I => \N__12255\
        );

    \I__2234\ : InMux
    port map (
            O => \N__12260\,
            I => \N__12252\
        );

    \I__2233\ : Span4Mux_v
    port map (
            O => \N__12255\,
            I => \N__12245\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__12252\,
            I => \N__12245\
        );

    \I__2231\ : InMux
    port map (
            O => \N__12251\,
            I => \N__12240\
        );

    \I__2230\ : InMux
    port map (
            O => \N__12250\,
            I => \N__12240\
        );

    \I__2229\ : Odrv4
    port map (
            O => \N__12245\,
            I => fifo_write_cmd
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__12240\,
            I => fifo_write_cmd
        );

    \I__2227\ : InMux
    port map (
            O => \N__12235\,
            I => \N__12230\
        );

    \I__2226\ : InMux
    port map (
            O => \N__12234\,
            I => \N__12225\
        );

    \I__2225\ : InMux
    port map (
            O => \N__12233\,
            I => \N__12225\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__12230\,
            I => wr_addr_r_2
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__12225\,
            I => wr_addr_r_2
        );

    \I__2222\ : InMux
    port map (
            O => \N__12220\,
            I => \N__12216\
        );

    \I__2221\ : InMux
    port map (
            O => \N__12219\,
            I => \N__12213\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__12216\,
            I => \N__12208\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__12213\,
            I => \N__12208\
        );

    \I__2218\ : Odrv4
    port map (
            O => \N__12208\,
            I => rd_addr_p1_w_1
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__12205\,
            I => \N__12201\
        );

    \I__2216\ : InMux
    port map (
            O => \N__12204\,
            I => \N__12198\
        );

    \I__2215\ : InMux
    port map (
            O => \N__12201\,
            I => \N__12195\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__12198\,
            I => rd_addr_p1_w_2
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__12195\,
            I => rd_addr_p1_w_2
        );

    \I__2212\ : CascadeMux
    port map (
            O => \N__12190\,
            I => \N__12183\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__12189\,
            I => \N__12178\
        );

    \I__2210\ : CascadeMux
    port map (
            O => \N__12188\,
            I => \N__12175\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__12187\,
            I => \N__12172\
        );

    \I__2208\ : InMux
    port map (
            O => \N__12186\,
            I => \N__12155\
        );

    \I__2207\ : InMux
    port map (
            O => \N__12183\,
            I => \N__12145\
        );

    \I__2206\ : InMux
    port map (
            O => \N__12182\,
            I => \N__12140\
        );

    \I__2205\ : InMux
    port map (
            O => \N__12181\,
            I => \N__12140\
        );

    \I__2204\ : InMux
    port map (
            O => \N__12178\,
            I => \N__12137\
        );

    \I__2203\ : InMux
    port map (
            O => \N__12175\,
            I => \N__12132\
        );

    \I__2202\ : InMux
    port map (
            O => \N__12172\,
            I => \N__12132\
        );

    \I__2201\ : InMux
    port map (
            O => \N__12171\,
            I => \N__12129\
        );

    \I__2200\ : InMux
    port map (
            O => \N__12170\,
            I => \N__12122\
        );

    \I__2199\ : InMux
    port map (
            O => \N__12169\,
            I => \N__12122\
        );

    \I__2198\ : InMux
    port map (
            O => \N__12168\,
            I => \N__12122\
        );

    \I__2197\ : InMux
    port map (
            O => \N__12167\,
            I => \N__12116\
        );

    \I__2196\ : InMux
    port map (
            O => \N__12166\,
            I => \N__12116\
        );

    \I__2195\ : InMux
    port map (
            O => \N__12165\,
            I => \N__12109\
        );

    \I__2194\ : InMux
    port map (
            O => \N__12164\,
            I => \N__12109\
        );

    \I__2193\ : InMux
    port map (
            O => \N__12163\,
            I => \N__12109\
        );

    \I__2192\ : InMux
    port map (
            O => \N__12162\,
            I => \N__12094\
        );

    \I__2191\ : InMux
    port map (
            O => \N__12161\,
            I => \N__12094\
        );

    \I__2190\ : InMux
    port map (
            O => \N__12160\,
            I => \N__12094\
        );

    \I__2189\ : InMux
    port map (
            O => \N__12159\,
            I => \N__12094\
        );

    \I__2188\ : InMux
    port map (
            O => \N__12158\,
            I => \N__12094\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__12155\,
            I => \N__12091\
        );

    \I__2186\ : InMux
    port map (
            O => \N__12154\,
            I => \N__12079\
        );

    \I__2185\ : InMux
    port map (
            O => \N__12153\,
            I => \N__12079\
        );

    \I__2184\ : InMux
    port map (
            O => \N__12152\,
            I => \N__12079\
        );

    \I__2183\ : InMux
    port map (
            O => \N__12151\,
            I => \N__12079\
        );

    \I__2182\ : InMux
    port map (
            O => \N__12150\,
            I => \N__12079\
        );

    \I__2181\ : InMux
    port map (
            O => \N__12149\,
            I => \N__12074\
        );

    \I__2180\ : InMux
    port map (
            O => \N__12148\,
            I => \N__12074\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__12145\,
            I => \N__12071\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__12140\,
            I => \N__12068\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__12137\,
            I => \N__12063\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__12132\,
            I => \N__12063\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__12129\,
            I => \N__12058\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__12122\,
            I => \N__12058\
        );

    \I__2173\ : CascadeMux
    port map (
            O => \N__12121\,
            I => \N__12054\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__12116\,
            I => \N__12049\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__12109\,
            I => \N__12049\
        );

    \I__2170\ : InMux
    port map (
            O => \N__12108\,
            I => \N__12040\
        );

    \I__2169\ : InMux
    port map (
            O => \N__12107\,
            I => \N__12040\
        );

    \I__2168\ : InMux
    port map (
            O => \N__12106\,
            I => \N__12040\
        );

    \I__2167\ : InMux
    port map (
            O => \N__12105\,
            I => \N__12040\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__12094\,
            I => \N__12035\
        );

    \I__2165\ : Span4Mux_v
    port map (
            O => \N__12091\,
            I => \N__12035\
        );

    \I__2164\ : CascadeMux
    port map (
            O => \N__12090\,
            I => \N__12031\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__12079\,
            I => \N__12026\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__12074\,
            I => \N__12026\
        );

    \I__2161\ : Span4Mux_v
    port map (
            O => \N__12071\,
            I => \N__12021\
        );

    \I__2160\ : Span4Mux_h
    port map (
            O => \N__12068\,
            I => \N__12021\
        );

    \I__2159\ : Span4Mux_v
    port map (
            O => \N__12063\,
            I => \N__12016\
        );

    \I__2158\ : Span4Mux_h
    port map (
            O => \N__12058\,
            I => \N__12016\
        );

    \I__2157\ : InMux
    port map (
            O => \N__12057\,
            I => \N__12011\
        );

    \I__2156\ : InMux
    port map (
            O => \N__12054\,
            I => \N__12008\
        );

    \I__2155\ : Span4Mux_v
    port map (
            O => \N__12049\,
            I => \N__12005\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__12040\,
            I => \N__12000\
        );

    \I__2153\ : Sp12to4
    port map (
            O => \N__12035\,
            I => \N__12000\
        );

    \I__2152\ : InMux
    port map (
            O => \N__12034\,
            I => \N__11995\
        );

    \I__2151\ : InMux
    port map (
            O => \N__12031\,
            I => \N__11995\
        );

    \I__2150\ : Span4Mux_h
    port map (
            O => \N__12026\,
            I => \N__11990\
        );

    \I__2149\ : Span4Mux_h
    port map (
            O => \N__12021\,
            I => \N__11990\
        );

    \I__2148\ : Span4Mux_h
    port map (
            O => \N__12016\,
            I => \N__11987\
        );

    \I__2147\ : InMux
    port map (
            O => \N__12015\,
            I => \N__11982\
        );

    \I__2146\ : InMux
    port map (
            O => \N__12014\,
            I => \N__11982\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__12011\,
            I => wr_addr_r_1
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__12008\,
            I => wr_addr_r_1
        );

    \I__2143\ : Odrv4
    port map (
            O => \N__12005\,
            I => wr_addr_r_1
        );

    \I__2142\ : Odrv12
    port map (
            O => \N__12000\,
            I => wr_addr_r_1
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__11995\,
            I => wr_addr_r_1
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__11990\,
            I => wr_addr_r_1
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__11987\,
            I => wr_addr_r_1
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__11982\,
            I => wr_addr_r_1
        );

    \I__2137\ : CascadeMux
    port map (
            O => \N__11965\,
            I => \n5474_cascade_\
        );

    \I__2136\ : InMux
    port map (
            O => \N__11962\,
            I => \N__11959\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__11959\,
            I => n24_adj_674
        );

    \I__2134\ : InMux
    port map (
            O => \N__11956\,
            I => \N__11946\
        );

    \I__2133\ : InMux
    port map (
            O => \N__11955\,
            I => \N__11946\
        );

    \I__2132\ : InMux
    port map (
            O => \N__11954\,
            I => \N__11937\
        );

    \I__2131\ : InMux
    port map (
            O => \N__11953\,
            I => \N__11937\
        );

    \I__2130\ : InMux
    port map (
            O => \N__11952\,
            I => \N__11937\
        );

    \I__2129\ : InMux
    port map (
            O => \N__11951\,
            I => \N__11933\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__11946\,
            I => \N__11930\
        );

    \I__2127\ : InMux
    port map (
            O => \N__11945\,
            I => \N__11925\
        );

    \I__2126\ : InMux
    port map (
            O => \N__11944\,
            I => \N__11925\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__11937\,
            I => \N__11922\
        );

    \I__2124\ : InMux
    port map (
            O => \N__11936\,
            I => \N__11919\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__11933\,
            I => wr_addr_r_0
        );

    \I__2122\ : Odrv12
    port map (
            O => \N__11930\,
            I => wr_addr_r_0
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__11925\,
            I => wr_addr_r_0
        );

    \I__2120\ : Odrv4
    port map (
            O => \N__11922\,
            I => wr_addr_r_0
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__11919\,
            I => wr_addr_r_0
        );

    \I__2118\ : InMux
    port map (
            O => \N__11908\,
            I => \N__11905\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__11905\,
            I => n4_adj_675
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__11902\,
            I => \N__11896\
        );

    \I__2115\ : InMux
    port map (
            O => \N__11901\,
            I => \N__11891\
        );

    \I__2114\ : InMux
    port map (
            O => \N__11900\,
            I => \N__11888\
        );

    \I__2113\ : InMux
    port map (
            O => \N__11899\,
            I => \N__11885\
        );

    \I__2112\ : InMux
    port map (
            O => \N__11896\,
            I => \N__11880\
        );

    \I__2111\ : InMux
    port map (
            O => \N__11895\,
            I => \N__11880\
        );

    \I__2110\ : CascadeMux
    port map (
            O => \N__11894\,
            I => \N__11877\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__11891\,
            I => \N__11873\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__11888\,
            I => \N__11870\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__11885\,
            I => \N__11865\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__11880\,
            I => \N__11865\
        );

    \I__2105\ : InMux
    port map (
            O => \N__11877\,
            I => \N__11860\
        );

    \I__2104\ : InMux
    port map (
            O => \N__11876\,
            I => \N__11860\
        );

    \I__2103\ : Span4Mux_v
    port map (
            O => \N__11873\,
            I => \N__11857\
        );

    \I__2102\ : Span4Mux_v
    port map (
            O => \N__11870\,
            I => \N__11850\
        );

    \I__2101\ : Span4Mux_h
    port map (
            O => \N__11865\,
            I => \N__11850\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__11860\,
            I => \N__11850\
        );

    \I__2099\ : Span4Mux_h
    port map (
            O => \N__11857\,
            I => \N__11846\
        );

    \I__2098\ : Span4Mux_v
    port map (
            O => \N__11850\,
            I => \N__11843\
        );

    \I__2097\ : InMux
    port map (
            O => \N__11849\,
            I => \N__11840\
        );

    \I__2096\ : Odrv4
    port map (
            O => \N__11846\,
            I => n2545
        );

    \I__2095\ : Odrv4
    port map (
            O => \N__11843\,
            I => n2545
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__11840\,
            I => n2545
        );

    \I__2093\ : CascadeMux
    port map (
            O => \N__11833\,
            I => \N__11830\
        );

    \I__2092\ : InMux
    port map (
            O => \N__11830\,
            I => \N__11827\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__11827\,
            I => \tx_fifo.lscc_fifo_inst.rd_fifo_en_prev_r\
        );

    \I__2090\ : CascadeMux
    port map (
            O => \N__11824\,
            I => \pc_rx.n5478_cascade_\
        );

    \I__2089\ : InMux
    port map (
            O => \N__11821\,
            I => \N__11818\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__11818\,
            I => \pc_rx.n6\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__11815\,
            I => \pc_rx.n5488_cascade_\
        );

    \I__2086\ : InMux
    port map (
            O => \N__11812\,
            I => \N__11806\
        );

    \I__2085\ : InMux
    port map (
            O => \N__11811\,
            I => \N__11806\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__11806\,
            I => \N__11802\
        );

    \I__2083\ : InMux
    port map (
            O => \N__11805\,
            I => \N__11799\
        );

    \I__2082\ : Odrv4
    port map (
            O => \N__11802\,
            I => \pc_rx.r_SM_Main_2_N_252_0\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__11799\,
            I => \pc_rx.r_SM_Main_2_N_252_0\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__11794\,
            I => \pc_rx.r_SM_Main_2_N_252_0_cascade_\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__11791\,
            I => \N__11788\
        );

    \I__2078\ : InMux
    port map (
            O => \N__11788\,
            I => \N__11785\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__11785\,
            I => \pc_rx.n6_adj_635\
        );

    \I__2076\ : CascadeMux
    port map (
            O => \N__11782\,
            I => \N__11779\
        );

    \I__2075\ : InMux
    port map (
            O => \N__11779\,
            I => \N__11776\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__11776\,
            I => \N__11773\
        );

    \I__2073\ : Span4Mux_h
    port map (
            O => \N__11773\,
            I => \N__11769\
        );

    \I__2072\ : InMux
    port map (
            O => \N__11772\,
            I => \N__11766\
        );

    \I__2071\ : Span4Mux_v
    port map (
            O => \N__11769\,
            I => \N__11762\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__11766\,
            I => \N__11759\
        );

    \I__2069\ : InMux
    port map (
            O => \N__11765\,
            I => \N__11756\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__11762\,
            I => tx_data_byte_7
        );

    \I__2067\ : Odrv4
    port map (
            O => \N__11759\,
            I => tx_data_byte_7
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__11756\,
            I => tx_data_byte_7
        );

    \I__2065\ : InMux
    port map (
            O => \N__11749\,
            I => \N__11745\
        );

    \I__2064\ : InMux
    port map (
            O => \N__11748\,
            I => \N__11742\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__11745\,
            I => tx_addr_byte_7
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__11742\,
            I => tx_addr_byte_7
        );

    \I__2061\ : InMux
    port map (
            O => \N__11737\,
            I => \N__11730\
        );

    \I__2060\ : InMux
    port map (
            O => \N__11736\,
            I => \N__11727\
        );

    \I__2059\ : InMux
    port map (
            O => \N__11735\,
            I => \N__11718\
        );

    \I__2058\ : InMux
    port map (
            O => \N__11734\,
            I => \N__11711\
        );

    \I__2057\ : InMux
    port map (
            O => \N__11733\,
            I => \N__11711\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__11730\,
            I => \N__11706\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__11727\,
            I => \N__11706\
        );

    \I__2054\ : InMux
    port map (
            O => \N__11726\,
            I => \N__11703\
        );

    \I__2053\ : InMux
    port map (
            O => \N__11725\,
            I => \N__11698\
        );

    \I__2052\ : InMux
    port map (
            O => \N__11724\,
            I => \N__11698\
        );

    \I__2051\ : InMux
    port map (
            O => \N__11723\,
            I => \N__11691\
        );

    \I__2050\ : InMux
    port map (
            O => \N__11722\,
            I => \N__11691\
        );

    \I__2049\ : InMux
    port map (
            O => \N__11721\,
            I => \N__11691\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__11718\,
            I => \N__11688\
        );

    \I__2047\ : InMux
    port map (
            O => \N__11717\,
            I => \N__11685\
        );

    \I__2046\ : InMux
    port map (
            O => \N__11716\,
            I => \N__11682\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__11711\,
            I => state_reg_0
        );

    \I__2044\ : Odrv4
    port map (
            O => \N__11706\,
            I => state_reg_0
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__11703\,
            I => state_reg_0
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__11698\,
            I => state_reg_0
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__11691\,
            I => state_reg_0
        );

    \I__2040\ : Odrv12
    port map (
            O => \N__11688\,
            I => state_reg_0
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__11685\,
            I => state_reg_0
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__11682\,
            I => state_reg_0
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__11665\,
            I => \N__11662\
        );

    \I__2036\ : InMux
    port map (
            O => \N__11662\,
            I => \N__11659\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__11659\,
            I => \N__11656\
        );

    \I__2034\ : Span4Mux_h
    port map (
            O => \N__11656\,
            I => \N__11652\
        );

    \I__2033\ : InMux
    port map (
            O => \N__11655\,
            I => \N__11649\
        );

    \I__2032\ : Odrv4
    port map (
            O => \N__11652\,
            I => tx_addr_byte_2
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__11649\,
            I => tx_addr_byte_2
        );

    \I__2030\ : InMux
    port map (
            O => \N__11644\,
            I => \N__11641\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__11641\,
            I => wr_addr_p1_w_2
        );

    \I__2028\ : CascadeMux
    port map (
            O => \N__11638\,
            I => \wr_addr_p1_w_2_cascade_\
        );

    \I__2027\ : InMux
    port map (
            O => \N__11635\,
            I => \N__11630\
        );

    \I__2026\ : InMux
    port map (
            O => \N__11634\,
            I => \N__11625\
        );

    \I__2025\ : InMux
    port map (
            O => \N__11633\,
            I => \N__11625\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__11630\,
            I => wr_fifo_en_w
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__11625\,
            I => wr_fifo_en_w
        );

    \I__2022\ : InMux
    port map (
            O => \N__11620\,
            I => \N__11617\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__11617\,
            I => \N__11614\
        );

    \I__2020\ : Span12Mux_v
    port map (
            O => \N__11614\,
            I => \N__11610\
        );

    \I__2019\ : InMux
    port map (
            O => \N__11613\,
            I => \N__11607\
        );

    \I__2018\ : Odrv12
    port map (
            O => \N__11610\,
            I => tx_addr_byte_5
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__11607\,
            I => tx_addr_byte_5
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__11602\,
            I => \N__11598\
        );

    \I__2015\ : InMux
    port map (
            O => \N__11601\,
            I => \N__11593\
        );

    \I__2014\ : InMux
    port map (
            O => \N__11598\,
            I => \N__11593\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__11593\,
            I => pc_data_rx_1
        );

    \I__2012\ : InMux
    port map (
            O => \N__11590\,
            I => \N__11587\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__11587\,
            I => \N__11582\
        );

    \I__2010\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11577\
        );

    \I__2009\ : InMux
    port map (
            O => \N__11585\,
            I => \N__11577\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__11582\,
            I => tx_data_byte_1
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__11577\,
            I => tx_data_byte_1
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__11572\,
            I => \pc_rx.n5452_cascade_\
        );

    \I__2005\ : InMux
    port map (
            O => \N__11569\,
            I => \N__11566\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__11566\,
            I => \N__11563\
        );

    \I__2003\ : Span4Mux_v
    port map (
            O => \N__11563\,
            I => \N__11560\
        );

    \I__2002\ : Sp12to4
    port map (
            O => \N__11560\,
            I => \N__11557\
        );

    \I__2001\ : Span12Mux_h
    port map (
            O => \N__11557\,
            I => \N__11554\
        );

    \I__2000\ : Odrv12
    port map (
            O => \N__11554\,
            I => \FIFO_D27_c_27\
        );

    \I__1999\ : IoInMux
    port map (
            O => \N__11551\,
            I => \N__11548\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__11548\,
            I => \N__11545\
        );

    \I__1997\ : Span4Mux_s1_v
    port map (
            O => \N__11545\,
            I => \N__11542\
        );

    \I__1996\ : Span4Mux_v
    port map (
            O => \N__11542\,
            I => \N__11539\
        );

    \I__1995\ : Span4Mux_v
    port map (
            O => \N__11539\,
            I => \N__11536\
        );

    \I__1994\ : Odrv4
    port map (
            O => \N__11536\,
            I => \DATA27_c_27\
        );

    \I__1993\ : InMux
    port map (
            O => \N__11533\,
            I => \N__11530\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__11530\,
            I => \N__11527\
        );

    \I__1991\ : Span4Mux_v
    port map (
            O => \N__11527\,
            I => \N__11524\
        );

    \I__1990\ : Sp12to4
    port map (
            O => \N__11524\,
            I => \N__11521\
        );

    \I__1989\ : Span12Mux_v
    port map (
            O => \N__11521\,
            I => \N__11518\
        );

    \I__1988\ : Span12Mux_h
    port map (
            O => \N__11518\,
            I => \N__11515\
        );

    \I__1987\ : Odrv12
    port map (
            O => \N__11515\,
            I => \FIFO_D20_c_20\
        );

    \I__1986\ : IoInMux
    port map (
            O => \N__11512\,
            I => \N__11509\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__11509\,
            I => \N__11506\
        );

    \I__1984\ : IoSpan4Mux
    port map (
            O => \N__11506\,
            I => \N__11503\
        );

    \I__1983\ : IoSpan4Mux
    port map (
            O => \N__11503\,
            I => \N__11500\
        );

    \I__1982\ : Span4Mux_s3_v
    port map (
            O => \N__11500\,
            I => \N__11497\
        );

    \I__1981\ : Sp12to4
    port map (
            O => \N__11497\,
            I => \N__11494\
        );

    \I__1980\ : Span12Mux_s11_v
    port map (
            O => \N__11494\,
            I => \N__11491\
        );

    \I__1979\ : Odrv12
    port map (
            O => \N__11491\,
            I => \DATA20_c_20\
        );

    \I__1978\ : InMux
    port map (
            O => \N__11488\,
            I => \N__11485\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__11485\,
            I => \N__11482\
        );

    \I__1976\ : Span4Mux_v
    port map (
            O => \N__11482\,
            I => \N__11479\
        );

    \I__1975\ : Sp12to4
    port map (
            O => \N__11479\,
            I => \N__11476\
        );

    \I__1974\ : Span12Mux_h
    port map (
            O => \N__11476\,
            I => \N__11473\
        );

    \I__1973\ : Span12Mux_v
    port map (
            O => \N__11473\,
            I => \N__11470\
        );

    \I__1972\ : Odrv12
    port map (
            O => \N__11470\,
            I => \FIFO_D13_c_13\
        );

    \I__1971\ : IoInMux
    port map (
            O => \N__11467\,
            I => \N__11464\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__11464\,
            I => \N__11461\
        );

    \I__1969\ : Span12Mux_s5_h
    port map (
            O => \N__11461\,
            I => \N__11458\
        );

    \I__1968\ : Span12Mux_h
    port map (
            O => \N__11458\,
            I => \N__11455\
        );

    \I__1967\ : Odrv12
    port map (
            O => \N__11455\,
            I => \DATA13_c_13\
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__11452\,
            I => \N__11449\
        );

    \I__1965\ : InMux
    port map (
            O => \N__11449\,
            I => \N__11446\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__11446\,
            I => \N__11443\
        );

    \I__1963\ : Span4Mux_v
    port map (
            O => \N__11443\,
            I => \N__11439\
        );

    \I__1962\ : InMux
    port map (
            O => \N__11442\,
            I => \N__11436\
        );

    \I__1961\ : Odrv4
    port map (
            O => \N__11439\,
            I => tx_addr_byte_4
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__11436\,
            I => tx_addr_byte_4
        );

    \I__1959\ : InMux
    port map (
            O => \N__11431\,
            I => \N__11428\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__11428\,
            I => \pc_rx.n5450\
        );

    \I__1957\ : InMux
    port map (
            O => \N__11425\,
            I => \N__11422\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__11422\,
            I => \pc_rx.n1\
        );

    \I__1955\ : InMux
    port map (
            O => \N__11419\,
            I => \N__11416\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__11416\,
            I => \N__11413\
        );

    \I__1953\ : Span4Mux_v
    port map (
            O => \N__11413\,
            I => \N__11409\
        );

    \I__1952\ : InMux
    port map (
            O => \N__11412\,
            I => \N__11406\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__11409\,
            I => tx_addr_byte_1
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__11406\,
            I => tx_addr_byte_1
        );

    \I__1949\ : IoInMux
    port map (
            O => \N__11401\,
            I => \N__11398\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__11398\,
            I => \N__11395\
        );

    \I__1947\ : IoSpan4Mux
    port map (
            O => \N__11395\,
            I => \N__11392\
        );

    \I__1946\ : Span4Mux_s2_v
    port map (
            O => \N__11392\,
            I => \N__11389\
        );

    \I__1945\ : Span4Mux_h
    port map (
            O => \N__11389\,
            I => \N__11386\
        );

    \I__1944\ : Sp12to4
    port map (
            O => \N__11386\,
            I => \N__11382\
        );

    \I__1943\ : InMux
    port map (
            O => \N__11385\,
            I => \N__11379\
        );

    \I__1942\ : Span12Mux_v
    port map (
            O => \N__11382\,
            I => \N__11376\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__11379\,
            I => \N__11373\
        );

    \I__1940\ : Odrv12
    port map (
            O => \N__11376\,
            I => \RESET_c\
        );

    \I__1939\ : Odrv4
    port map (
            O => \N__11373\,
            I => \RESET_c\
        );

    \I__1938\ : CascadeMux
    port map (
            O => \N__11368\,
            I => \n15_adj_673_cascade_\
        );

    \I__1937\ : InMux
    port map (
            O => \N__11365\,
            I => \N__11362\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__11362\,
            I => n4892
        );

    \I__1935\ : InMux
    port map (
            O => \N__11359\,
            I => \N__11350\
        );

    \I__1934\ : InMux
    port map (
            O => \N__11358\,
            I => \N__11350\
        );

    \I__1933\ : InMux
    port map (
            O => \N__11357\,
            I => \N__11350\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__11350\,
            I => \tx_fifo.lscc_fifo_inst.rd_addr_r_2\
        );

    \I__1931\ : InMux
    port map (
            O => \N__11347\,
            I => \N__11341\
        );

    \I__1930\ : InMux
    port map (
            O => \N__11346\,
            I => \N__11341\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__11341\,
            I => n1
        );

    \I__1928\ : CEMux
    port map (
            O => \N__11338\,
            I => \N__11335\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__11335\,
            I => \N__11331\
        );

    \I__1926\ : CEMux
    port map (
            O => \N__11334\,
            I => \N__11327\
        );

    \I__1925\ : Span4Mux_h
    port map (
            O => \N__11331\,
            I => \N__11324\
        );

    \I__1924\ : CEMux
    port map (
            O => \N__11330\,
            I => \N__11321\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__11327\,
            I => \N__11317\
        );

    \I__1922\ : Span4Mux_v
    port map (
            O => \N__11324\,
            I => \N__11312\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__11321\,
            I => \N__11312\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__11320\,
            I => \N__11309\
        );

    \I__1919\ : Span4Mux_h
    port map (
            O => \N__11317\,
            I => \N__11306\
        );

    \I__1918\ : Span4Mux_h
    port map (
            O => \N__11312\,
            I => \N__11303\
        );

    \I__1917\ : InMux
    port map (
            O => \N__11309\,
            I => \N__11300\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__11306\,
            I => \tx_fifo.lscc_fifo_inst.rd_fifo_en_w\
        );

    \I__1915\ : Odrv4
    port map (
            O => \N__11303\,
            I => \tx_fifo.lscc_fifo_inst.rd_fifo_en_w\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__11300\,
            I => \tx_fifo.lscc_fifo_inst.rd_fifo_en_w\
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__11293\,
            I => \tx_fifo.lscc_fifo_inst.rd_fifo_en_w_cascade_\
        );

    \I__1912\ : CascadeMux
    port map (
            O => \N__11290\,
            I => \N__11287\
        );

    \I__1911\ : InMux
    port map (
            O => \N__11287\,
            I => \N__11284\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__11284\,
            I => \N__11281\
        );

    \I__1909\ : Span4Mux_h
    port map (
            O => \N__11281\,
            I => \N__11278\
        );

    \I__1908\ : Odrv4
    port map (
            O => \N__11278\,
            I => \mem_LUT_data_raw_r_7\
        );

    \I__1907\ : InMux
    port map (
            O => \N__11275\,
            I => \N__11272\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__11272\,
            I => \N__11269\
        );

    \I__1905\ : Span4Mux_h
    port map (
            O => \N__11269\,
            I => \N__11266\
        );

    \I__1904\ : Span4Mux_v
    port map (
            O => \N__11266\,
            I => \N__11262\
        );

    \I__1903\ : InMux
    port map (
            O => \N__11265\,
            I => \N__11259\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__11262\,
            I => fifo_temp_output_7
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__11259\,
            I => fifo_temp_output_7
        );

    \I__1900\ : CascadeMux
    port map (
            O => \N__11254\,
            I => \N__11251\
        );

    \I__1899\ : InMux
    port map (
            O => \N__11251\,
            I => \N__11244\
        );

    \I__1898\ : InMux
    port map (
            O => \N__11250\,
            I => \N__11237\
        );

    \I__1897\ : InMux
    port map (
            O => \N__11249\,
            I => \N__11237\
        );

    \I__1896\ : InMux
    port map (
            O => \N__11248\,
            I => \N__11237\
        );

    \I__1895\ : InMux
    port map (
            O => \N__11247\,
            I => \N__11233\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__11244\,
            I => \N__11228\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__11237\,
            I => \N__11228\
        );

    \I__1892\ : InMux
    port map (
            O => \N__11236\,
            I => \N__11225\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__11233\,
            I => is_tx_fifo_full_flag
        );

    \I__1890\ : Odrv12
    port map (
            O => \N__11228\,
            I => is_tx_fifo_full_flag
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__11225\,
            I => is_tx_fifo_full_flag
        );

    \I__1888\ : InMux
    port map (
            O => \N__11218\,
            I => \N__11215\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__11215\,
            I => \N__11212\
        );

    \I__1886\ : Odrv12
    port map (
            O => \N__11212\,
            I => tx_shift_reg_11
        );

    \I__1885\ : InMux
    port map (
            O => \N__11209\,
            I => \N__11206\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__11206\,
            I => tx_shift_reg_2
        );

    \I__1883\ : InMux
    port map (
            O => \N__11203\,
            I => \N__11200\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__11200\,
            I => tx_shift_reg_12
        );

    \I__1881\ : InMux
    port map (
            O => \N__11197\,
            I => \N__11194\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__11194\,
            I => tx_shift_reg_13
        );

    \I__1879\ : InMux
    port map (
            O => \N__11191\,
            I => \N__11188\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__11188\,
            I => tx_shift_reg_14
        );

    \I__1877\ : InMux
    port map (
            O => \N__11185\,
            I => \N__11182\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__11182\,
            I => \N__11173\
        );

    \I__1875\ : InMux
    port map (
            O => \N__11181\,
            I => \N__11170\
        );

    \I__1874\ : InMux
    port map (
            O => \N__11180\,
            I => \N__11157\
        );

    \I__1873\ : InMux
    port map (
            O => \N__11179\,
            I => \N__11157\
        );

    \I__1872\ : InMux
    port map (
            O => \N__11178\,
            I => \N__11157\
        );

    \I__1871\ : InMux
    port map (
            O => \N__11177\,
            I => \N__11157\
        );

    \I__1870\ : InMux
    port map (
            O => \N__11176\,
            I => \N__11157\
        );

    \I__1869\ : Span4Mux_v
    port map (
            O => \N__11173\,
            I => \N__11152\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__11170\,
            I => \N__11152\
        );

    \I__1867\ : InMux
    port map (
            O => \N__11169\,
            I => \N__11147\
        );

    \I__1866\ : InMux
    port map (
            O => \N__11168\,
            I => \N__11147\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__11157\,
            I => \N__11140\
        );

    \I__1864\ : Span4Mux_v
    port map (
            O => \N__11152\,
            I => \N__11140\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__11147\,
            I => \N__11140\
        );

    \I__1862\ : Span4Mux_h
    port map (
            O => \N__11140\,
            I => \N__11123\
        );

    \I__1861\ : InMux
    port map (
            O => \N__11139\,
            I => \N__11110\
        );

    \I__1860\ : InMux
    port map (
            O => \N__11138\,
            I => \N__11110\
        );

    \I__1859\ : InMux
    port map (
            O => \N__11137\,
            I => \N__11110\
        );

    \I__1858\ : InMux
    port map (
            O => \N__11136\,
            I => \N__11110\
        );

    \I__1857\ : InMux
    port map (
            O => \N__11135\,
            I => \N__11110\
        );

    \I__1856\ : InMux
    port map (
            O => \N__11134\,
            I => \N__11110\
        );

    \I__1855\ : InMux
    port map (
            O => \N__11133\,
            I => \N__11095\
        );

    \I__1854\ : InMux
    port map (
            O => \N__11132\,
            I => \N__11095\
        );

    \I__1853\ : InMux
    port map (
            O => \N__11131\,
            I => \N__11095\
        );

    \I__1852\ : InMux
    port map (
            O => \N__11130\,
            I => \N__11095\
        );

    \I__1851\ : InMux
    port map (
            O => \N__11129\,
            I => \N__11095\
        );

    \I__1850\ : InMux
    port map (
            O => \N__11128\,
            I => \N__11095\
        );

    \I__1849\ : InMux
    port map (
            O => \N__11127\,
            I => \N__11095\
        );

    \I__1848\ : InMux
    port map (
            O => \N__11126\,
            I => \N__11092\
        );

    \I__1847\ : Odrv4
    port map (
            O => \N__11123\,
            I => n5462
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__11110\,
            I => n5462
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__11095\,
            I => n5462
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__11092\,
            I => n5462
        );

    \I__1843\ : CascadeMux
    port map (
            O => \N__11083\,
            I => \N__11072\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__11082\,
            I => \N__11069\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__11081\,
            I => \N__11065\
        );

    \I__1840\ : CascadeMux
    port map (
            O => \N__11080\,
            I => \N__11061\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__11079\,
            I => \N__11058\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__11078\,
            I => \N__11053\
        );

    \I__1837\ : InMux
    port map (
            O => \N__11077\,
            I => \N__11047\
        );

    \I__1836\ : InMux
    port map (
            O => \N__11076\,
            I => \N__11047\
        );

    \I__1835\ : InMux
    port map (
            O => \N__11075\,
            I => \N__11034\
        );

    \I__1834\ : InMux
    port map (
            O => \N__11072\,
            I => \N__11034\
        );

    \I__1833\ : InMux
    port map (
            O => \N__11069\,
            I => \N__11034\
        );

    \I__1832\ : InMux
    port map (
            O => \N__11068\,
            I => \N__11034\
        );

    \I__1831\ : InMux
    port map (
            O => \N__11065\,
            I => \N__11034\
        );

    \I__1830\ : InMux
    port map (
            O => \N__11064\,
            I => \N__11034\
        );

    \I__1829\ : InMux
    port map (
            O => \N__11061\,
            I => \N__11021\
        );

    \I__1828\ : InMux
    port map (
            O => \N__11058\,
            I => \N__11021\
        );

    \I__1827\ : InMux
    port map (
            O => \N__11057\,
            I => \N__11021\
        );

    \I__1826\ : InMux
    port map (
            O => \N__11056\,
            I => \N__11021\
        );

    \I__1825\ : InMux
    port map (
            O => \N__11053\,
            I => \N__11021\
        );

    \I__1824\ : InMux
    port map (
            O => \N__11052\,
            I => \N__11021\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__11047\,
            I => n2446
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__11034\,
            I => n2446
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__11021\,
            I => n2446
        );

    \I__1820\ : InMux
    port map (
            O => \N__11014\,
            I => \N__11011\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__11011\,
            I => tx_shift_reg_1
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__11008\,
            I => \N__11004\
        );

    \I__1817\ : InMux
    port map (
            O => \N__11007\,
            I => \N__11001\
        );

    \I__1816\ : InMux
    port map (
            O => \N__11004\,
            I => \N__10998\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__11001\,
            I => \N__10995\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__10998\,
            I => \N__10991\
        );

    \I__1813\ : Span4Mux_v
    port map (
            O => \N__10995\,
            I => \N__10988\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__10994\,
            I => \N__10985\
        );

    \I__1811\ : Span4Mux_v
    port map (
            O => \N__10991\,
            I => \N__10982\
        );

    \I__1810\ : Span4Mux_h
    port map (
            O => \N__10988\,
            I => \N__10979\
        );

    \I__1809\ : InMux
    port map (
            O => \N__10985\,
            I => \N__10976\
        );

    \I__1808\ : Odrv4
    port map (
            O => \N__10982\,
            I => tx_uart_active_flag
        );

    \I__1807\ : Odrv4
    port map (
            O => \N__10979\,
            I => tx_uart_active_flag
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__10976\,
            I => tx_uart_active_flag
        );

    \I__1805\ : CascadeMux
    port map (
            O => \N__10969\,
            I => \n5454_cascade_\
        );

    \I__1804\ : InMux
    port map (
            O => \N__10966\,
            I => \N__10962\
        );

    \I__1803\ : InMux
    port map (
            O => \N__10965\,
            I => \N__10959\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__10962\,
            I => \pc_tx.r_Clock_Count_3\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__10959\,
            I => \pc_tx.r_Clock_Count_3\
        );

    \I__1800\ : InMux
    port map (
            O => \N__10954\,
            I => \pc_tx.n4867\
        );

    \I__1799\ : InMux
    port map (
            O => \N__10951\,
            I => \N__10947\
        );

    \I__1798\ : InMux
    port map (
            O => \N__10950\,
            I => \N__10944\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__10947\,
            I => \pc_tx.r_Clock_Count_4\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__10944\,
            I => \pc_tx.r_Clock_Count_4\
        );

    \I__1795\ : InMux
    port map (
            O => \N__10939\,
            I => \pc_tx.n4868\
        );

    \I__1794\ : InMux
    port map (
            O => \N__10936\,
            I => \N__10932\
        );

    \I__1793\ : InMux
    port map (
            O => \N__10935\,
            I => \N__10929\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__10932\,
            I => \pc_tx.r_Clock_Count_5\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__10929\,
            I => \pc_tx.r_Clock_Count_5\
        );

    \I__1790\ : InMux
    port map (
            O => \N__10924\,
            I => \pc_tx.n4869\
        );

    \I__1789\ : InMux
    port map (
            O => \N__10921\,
            I => \N__10917\
        );

    \I__1788\ : InMux
    port map (
            O => \N__10920\,
            I => \N__10914\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__10917\,
            I => \pc_tx.r_Clock_Count_6\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__10914\,
            I => \pc_tx.r_Clock_Count_6\
        );

    \I__1785\ : InMux
    port map (
            O => \N__10909\,
            I => \pc_tx.n4870\
        );

    \I__1784\ : InMux
    port map (
            O => \N__10906\,
            I => \N__10902\
        );

    \I__1783\ : InMux
    port map (
            O => \N__10905\,
            I => \N__10899\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__10902\,
            I => \pc_tx.r_Clock_Count_7\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__10899\,
            I => \pc_tx.r_Clock_Count_7\
        );

    \I__1780\ : InMux
    port map (
            O => \N__10894\,
            I => \pc_tx.n4871\
        );

    \I__1779\ : InMux
    port map (
            O => \N__10891\,
            I => \N__10887\
        );

    \I__1778\ : InMux
    port map (
            O => \N__10890\,
            I => \N__10884\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__10887\,
            I => \pc_tx.r_Clock_Count_8\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__10884\,
            I => \pc_tx.r_Clock_Count_8\
        );

    \I__1775\ : InMux
    port map (
            O => \N__10879\,
            I => \bfn_11_7_0_\
        );

    \I__1774\ : InMux
    port map (
            O => \N__10876\,
            I => \pc_tx.n4873\
        );

    \I__1773\ : InMux
    port map (
            O => \N__10873\,
            I => \N__10869\
        );

    \I__1772\ : InMux
    port map (
            O => \N__10872\,
            I => \N__10866\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__10869\,
            I => \pc_tx.r_Clock_Count_9\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__10866\,
            I => \pc_tx.r_Clock_Count_9\
        );

    \I__1769\ : SRMux
    port map (
            O => \N__10861\,
            I => \N__10858\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__10858\,
            I => \N__10854\
        );

    \I__1767\ : SRMux
    port map (
            O => \N__10857\,
            I => \N__10851\
        );

    \I__1766\ : Span4Mux_h
    port map (
            O => \N__10854\,
            I => \N__10846\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__10851\,
            I => \N__10846\
        );

    \I__1764\ : Odrv4
    port map (
            O => \N__10846\,
            I => \pc_tx.n2739\
        );

    \I__1763\ : IoInMux
    port map (
            O => \N__10843\,
            I => \N__10840\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__10840\,
            I => \N__10836\
        );

    \I__1761\ : IoInMux
    port map (
            O => \N__10839\,
            I => \N__10833\
        );

    \I__1760\ : Span4Mux_s2_v
    port map (
            O => \N__10836\,
            I => \N__10830\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__10833\,
            I => \N__10827\
        );

    \I__1758\ : Span4Mux_v
    port map (
            O => \N__10830\,
            I => \N__10824\
        );

    \I__1757\ : IoSpan4Mux
    port map (
            O => \N__10827\,
            I => \N__10821\
        );

    \I__1756\ : Span4Mux_v
    port map (
            O => \N__10824\,
            I => \N__10818\
        );

    \I__1755\ : Sp12to4
    port map (
            O => \N__10821\,
            I => \N__10815\
        );

    \I__1754\ : Sp12to4
    port map (
            O => \N__10818\,
            I => \N__10812\
        );

    \I__1753\ : Span12Mux_s9_v
    port map (
            O => \N__10815\,
            I => \N__10809\
        );

    \I__1752\ : Span12Mux_h
    port map (
            O => \N__10812\,
            I => \N__10804\
        );

    \I__1751\ : Span12Mux_h
    port map (
            O => \N__10809\,
            I => \N__10804\
        );

    \I__1750\ : Odrv12
    port map (
            O => \N__10804\,
            I => \DEBUG_9_c\
        );

    \I__1749\ : InMux
    port map (
            O => \N__10801\,
            I => \N__10798\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__10798\,
            I => \N__10795\
        );

    \I__1747\ : Span12Mux_h
    port map (
            O => \N__10795\,
            I => \N__10792\
        );

    \I__1746\ : Span12Mux_v
    port map (
            O => \N__10792\,
            I => \N__10789\
        );

    \I__1745\ : Odrv12
    port map (
            O => \N__10789\,
            I => \FIFO_D15_c_15\
        );

    \I__1744\ : IoInMux
    port map (
            O => \N__10786\,
            I => \N__10783\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__10783\,
            I => \N__10780\
        );

    \I__1742\ : IoSpan4Mux
    port map (
            O => \N__10780\,
            I => \N__10777\
        );

    \I__1741\ : Span4Mux_s2_h
    port map (
            O => \N__10777\,
            I => \N__10774\
        );

    \I__1740\ : Span4Mux_h
    port map (
            O => \N__10774\,
            I => \N__10771\
        );

    \I__1739\ : Sp12to4
    port map (
            O => \N__10771\,
            I => \N__10768\
        );

    \I__1738\ : Span12Mux_h
    port map (
            O => \N__10768\,
            I => \N__10765\
        );

    \I__1737\ : Odrv12
    port map (
            O => \N__10765\,
            I => \DATA15_c_15\
        );

    \I__1736\ : InMux
    port map (
            O => \N__10762\,
            I => \N__10756\
        );

    \I__1735\ : InMux
    port map (
            O => \N__10761\,
            I => \N__10756\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__10756\,
            I => \N__10753\
        );

    \I__1733\ : Span4Mux_v
    port map (
            O => \N__10753\,
            I => \N__10750\
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__10750\,
            I => spi_busy
        );

    \I__1731\ : InMux
    port map (
            O => \N__10747\,
            I => \N__10744\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__10744\,
            I => spi_busy_prev
        );

    \I__1729\ : CascadeMux
    port map (
            O => \N__10741\,
            I => \N__10736\
        );

    \I__1728\ : InMux
    port map (
            O => \N__10740\,
            I => \N__10730\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__10739\,
            I => \N__10725\
        );

    \I__1726\ : InMux
    port map (
            O => \N__10736\,
            I => \N__10718\
        );

    \I__1725\ : InMux
    port map (
            O => \N__10735\,
            I => \N__10711\
        );

    \I__1724\ : InMux
    port map (
            O => \N__10734\,
            I => \N__10711\
        );

    \I__1723\ : InMux
    port map (
            O => \N__10733\,
            I => \N__10711\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__10730\,
            I => \N__10708\
        );

    \I__1721\ : InMux
    port map (
            O => \N__10729\,
            I => \N__10705\
        );

    \I__1720\ : InMux
    port map (
            O => \N__10728\,
            I => \N__10702\
        );

    \I__1719\ : InMux
    port map (
            O => \N__10725\,
            I => \N__10693\
        );

    \I__1718\ : InMux
    port map (
            O => \N__10724\,
            I => \N__10693\
        );

    \I__1717\ : InMux
    port map (
            O => \N__10723\,
            I => \N__10688\
        );

    \I__1716\ : InMux
    port map (
            O => \N__10722\,
            I => \N__10688\
        );

    \I__1715\ : InMux
    port map (
            O => \N__10721\,
            I => \N__10685\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__10718\,
            I => \N__10674\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__10711\,
            I => \N__10674\
        );

    \I__1712\ : Span4Mux_h
    port map (
            O => \N__10708\,
            I => \N__10674\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__10705\,
            I => \N__10674\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__10702\,
            I => \N__10674\
        );

    \I__1709\ : InMux
    port map (
            O => \N__10701\,
            I => \N__10669\
        );

    \I__1708\ : InMux
    port map (
            O => \N__10700\,
            I => \N__10669\
        );

    \I__1707\ : InMux
    port map (
            O => \N__10699\,
            I => \N__10666\
        );

    \I__1706\ : InMux
    port map (
            O => \N__10698\,
            I => \N__10663\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__10693\,
            I => \N__10660\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__10688\,
            I => \N__10655\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__10685\,
            I => \N__10655\
        );

    \I__1702\ : Span4Mux_v
    port map (
            O => \N__10674\,
            I => \N__10650\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__10669\,
            I => \N__10650\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__10666\,
            I => \N__10645\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__10663\,
            I => \N__10645\
        );

    \I__1698\ : Span4Mux_v
    port map (
            O => \N__10660\,
            I => \N__10640\
        );

    \I__1697\ : Span4Mux_h
    port map (
            O => \N__10655\,
            I => \N__10640\
        );

    \I__1696\ : Span4Mux_h
    port map (
            O => \N__10650\,
            I => \N__10637\
        );

    \I__1695\ : Odrv12
    port map (
            O => \N__10645\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__10640\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__10637\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__1692\ : InMux
    port map (
            O => \N__10630\,
            I => \N__10627\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__10627\,
            I => spi_busy_falling_edge
        );

    \I__1690\ : CascadeMux
    port map (
            O => \N__10624\,
            I => \N__10618\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__10623\,
            I => \N__10609\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__10622\,
            I => \N__10606\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__10621\,
            I => \N__10601\
        );

    \I__1686\ : InMux
    port map (
            O => \N__10618\,
            I => \N__10596\
        );

    \I__1685\ : InMux
    port map (
            O => \N__10617\,
            I => \N__10593\
        );

    \I__1684\ : InMux
    port map (
            O => \N__10616\,
            I => \N__10582\
        );

    \I__1683\ : InMux
    port map (
            O => \N__10615\,
            I => \N__10582\
        );

    \I__1682\ : InMux
    port map (
            O => \N__10614\,
            I => \N__10582\
        );

    \I__1681\ : InMux
    port map (
            O => \N__10613\,
            I => \N__10582\
        );

    \I__1680\ : InMux
    port map (
            O => \N__10612\,
            I => \N__10582\
        );

    \I__1679\ : InMux
    port map (
            O => \N__10609\,
            I => \N__10573\
        );

    \I__1678\ : InMux
    port map (
            O => \N__10606\,
            I => \N__10573\
        );

    \I__1677\ : InMux
    port map (
            O => \N__10605\,
            I => \N__10573\
        );

    \I__1676\ : InMux
    port map (
            O => \N__10604\,
            I => \N__10573\
        );

    \I__1675\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10566\
        );

    \I__1674\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10566\
        );

    \I__1673\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10563\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__10596\,
            I => \N__10560\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__10593\,
            I => \N__10557\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__10582\,
            I => \N__10554\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__10573\,
            I => \N__10551\
        );

    \I__1668\ : InMux
    port map (
            O => \N__10572\,
            I => \N__10548\
        );

    \I__1667\ : InMux
    port map (
            O => \N__10571\,
            I => \N__10545\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__10566\,
            I => \N__10542\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__10563\,
            I => \N__10535\
        );

    \I__1664\ : Span4Mux_v
    port map (
            O => \N__10560\,
            I => \N__10535\
        );

    \I__1663\ : Span4Mux_v
    port map (
            O => \N__10557\,
            I => \N__10535\
        );

    \I__1662\ : Span4Mux_h
    port map (
            O => \N__10554\,
            I => \N__10532\
        );

    \I__1661\ : Span4Mux_v
    port map (
            O => \N__10551\,
            I => \N__10529\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__10548\,
            I => \N__10524\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__10545\,
            I => \N__10524\
        );

    \I__1658\ : Span4Mux_h
    port map (
            O => \N__10542\,
            I => \N__10521\
        );

    \I__1657\ : Span4Mux_h
    port map (
            O => \N__10535\,
            I => \N__10518\
        );

    \I__1656\ : Span4Mux_v
    port map (
            O => \N__10532\,
            I => \N__10515\
        );

    \I__1655\ : Span4Mux_h
    port map (
            O => \N__10529\,
            I => \N__10512\
        );

    \I__1654\ : Odrv12
    port map (
            O => \N__10524\,
            I => \tx_fifo.lscc_fifo_inst.n3\
        );

    \I__1653\ : Odrv4
    port map (
            O => \N__10521\,
            I => \tx_fifo.lscc_fifo_inst.n3\
        );

    \I__1652\ : Odrv4
    port map (
            O => \N__10518\,
            I => \tx_fifo.lscc_fifo_inst.n3\
        );

    \I__1651\ : Odrv4
    port map (
            O => \N__10515\,
            I => \tx_fifo.lscc_fifo_inst.n3\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__10512\,
            I => \tx_fifo.lscc_fifo_inst.n3\
        );

    \I__1649\ : InMux
    port map (
            O => \N__10501\,
            I => \N__10497\
        );

    \I__1648\ : InMux
    port map (
            O => \N__10500\,
            I => \N__10494\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__10497\,
            I => \pc_tx.r_Clock_Count_0\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__10494\,
            I => \pc_tx.r_Clock_Count_0\
        );

    \I__1645\ : InMux
    port map (
            O => \N__10489\,
            I => \bfn_11_6_0_\
        );

    \I__1644\ : InMux
    port map (
            O => \N__10486\,
            I => \N__10482\
        );

    \I__1643\ : InMux
    port map (
            O => \N__10485\,
            I => \N__10479\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__10482\,
            I => \pc_tx.r_Clock_Count_1\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__10479\,
            I => \pc_tx.r_Clock_Count_1\
        );

    \I__1640\ : InMux
    port map (
            O => \N__10474\,
            I => \pc_tx.n4865\
        );

    \I__1639\ : InMux
    port map (
            O => \N__10471\,
            I => \N__10467\
        );

    \I__1638\ : InMux
    port map (
            O => \N__10470\,
            I => \N__10464\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__10467\,
            I => \pc_tx.r_Clock_Count_2\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__10464\,
            I => \pc_tx.r_Clock_Count_2\
        );

    \I__1635\ : InMux
    port map (
            O => \N__10459\,
            I => \pc_tx.n4866\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__10456\,
            I => \N__10452\
        );

    \I__1633\ : InMux
    port map (
            O => \N__10455\,
            I => \N__10446\
        );

    \I__1632\ : InMux
    port map (
            O => \N__10452\,
            I => \N__10446\
        );

    \I__1631\ : InMux
    port map (
            O => \N__10451\,
            I => \N__10443\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__10446\,
            I => \reset_all_w_N_61\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__10443\,
            I => \reset_all_w_N_61\
        );

    \I__1628\ : InMux
    port map (
            O => \N__10438\,
            I => \N__10420\
        );

    \I__1627\ : InMux
    port map (
            O => \N__10437\,
            I => \N__10420\
        );

    \I__1626\ : InMux
    port map (
            O => \N__10436\,
            I => \N__10420\
        );

    \I__1625\ : InMux
    port map (
            O => \N__10435\,
            I => \N__10420\
        );

    \I__1624\ : InMux
    port map (
            O => \N__10434\,
            I => \N__10420\
        );

    \I__1623\ : InMux
    port map (
            O => \N__10433\,
            I => \N__10420\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__10420\,
            I => reset_clk_counter_0
        );

    \I__1621\ : CascadeMux
    port map (
            O => \N__10417\,
            I => \reset_all_w_N_61_cascade_\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__10414\,
            I => \N__10407\
        );

    \I__1619\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10404\
        );

    \I__1618\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10395\
        );

    \I__1617\ : InMux
    port map (
            O => \N__10411\,
            I => \N__10395\
        );

    \I__1616\ : InMux
    port map (
            O => \N__10410\,
            I => \N__10395\
        );

    \I__1615\ : InMux
    port map (
            O => \N__10407\,
            I => \N__10395\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__10404\,
            I => reset_clk_counter_1
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__10395\,
            I => reset_clk_counter_1
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__10390\,
            I => \n2_adj_670_cascade_\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__10387\,
            I => \N__10383\
        );

    \I__1610\ : InMux
    port map (
            O => \N__10386\,
            I => \N__10372\
        );

    \I__1609\ : InMux
    port map (
            O => \N__10383\,
            I => \N__10372\
        );

    \I__1608\ : InMux
    port map (
            O => \N__10382\,
            I => \N__10372\
        );

    \I__1607\ : InMux
    port map (
            O => \N__10381\,
            I => \N__10372\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__10372\,
            I => reset_clk_counter_2
        );

    \I__1605\ : InMux
    port map (
            O => \N__10369\,
            I => \N__10360\
        );

    \I__1604\ : InMux
    port map (
            O => \N__10368\,
            I => \N__10360\
        );

    \I__1603\ : InMux
    port map (
            O => \N__10367\,
            I => \N__10360\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__10360\,
            I => reset_clk_counter_3
        );

    \I__1601\ : InMux
    port map (
            O => \N__10357\,
            I => \N__10354\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__10354\,
            I => \N__10351\
        );

    \I__1599\ : Span4Mux_v
    port map (
            O => \N__10351\,
            I => \N__10348\
        );

    \I__1598\ : Span4Mux_h
    port map (
            O => \N__10348\,
            I => \N__10345\
        );

    \I__1597\ : Sp12to4
    port map (
            O => \N__10345\,
            I => \N__10342\
        );

    \I__1596\ : Odrv12
    port map (
            O => \N__10342\,
            I => \FIFO_D26_c_26\
        );

    \I__1595\ : IoInMux
    port map (
            O => \N__10339\,
            I => \N__10336\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__10336\,
            I => \N__10333\
        );

    \I__1593\ : Span12Mux_s2_v
    port map (
            O => \N__10333\,
            I => \N__10330\
        );

    \I__1592\ : Span12Mux_v
    port map (
            O => \N__10330\,
            I => \N__10327\
        );

    \I__1591\ : Odrv12
    port map (
            O => \N__10327\,
            I => \DATA26_c_26\
        );

    \I__1590\ : InMux
    port map (
            O => \N__10324\,
            I => \N__10321\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__10321\,
            I => tx_shift_reg_9
        );

    \I__1588\ : InMux
    port map (
            O => \N__10318\,
            I => \N__10315\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__10315\,
            I => tx_shift_reg_10
        );

    \I__1586\ : InMux
    port map (
            O => \N__10312\,
            I => \N__10309\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__10309\,
            I => tx_shift_reg_5
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__10306\,
            I => \n5462_cascade_\
        );

    \I__1583\ : InMux
    port map (
            O => \N__10303\,
            I => \N__10300\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__10300\,
            I => \N__10297\
        );

    \I__1581\ : Odrv4
    port map (
            O => \N__10297\,
            I => tx_shift_reg_6
        );

    \I__1580\ : InMux
    port map (
            O => \N__10294\,
            I => \N__10291\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__10291\,
            I => tx_shift_reg_7
        );

    \I__1578\ : InMux
    port map (
            O => \N__10288\,
            I => \N__10285\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__10285\,
            I => \N__10279\
        );

    \I__1576\ : InMux
    port map (
            O => \N__10284\,
            I => \N__10276\
        );

    \I__1575\ : InMux
    port map (
            O => \N__10283\,
            I => \N__10271\
        );

    \I__1574\ : InMux
    port map (
            O => \N__10282\,
            I => \N__10271\
        );

    \I__1573\ : Span4Mux_h
    port map (
            O => \N__10279\,
            I => \N__10268\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__10276\,
            I => \N__10263\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__10271\,
            I => \N__10263\
        );

    \I__1570\ : Span4Mux_v
    port map (
            O => \N__10268\,
            I => \N__10257\
        );

    \I__1569\ : Span4Mux_v
    port map (
            O => \N__10263\,
            I => \N__10257\
        );

    \I__1568\ : InMux
    port map (
            O => \N__10262\,
            I => \N__10254\
        );

    \I__1567\ : Odrv4
    port map (
            O => \N__10257\,
            I => rx_buf_byte_7
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__10254\,
            I => rx_buf_byte_7
        );

    \I__1565\ : InMux
    port map (
            O => \N__10249\,
            I => \N__10245\
        );

    \I__1564\ : InMux
    port map (
            O => \N__10248\,
            I => \N__10242\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__10245\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_7\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__10242\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_7\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__10237\,
            I => \N__10232\
        );

    \I__1560\ : CascadeMux
    port map (
            O => \N__10236\,
            I => \N__10229\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__10235\,
            I => \N__10226\
        );

    \I__1558\ : InMux
    port map (
            O => \N__10232\,
            I => \N__10221\
        );

    \I__1557\ : InMux
    port map (
            O => \N__10229\,
            I => \N__10221\
        );

    \I__1556\ : InMux
    port map (
            O => \N__10226\,
            I => \N__10218\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__10221\,
            I => \N__10214\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__10218\,
            I => \N__10211\
        );

    \I__1553\ : InMux
    port map (
            O => \N__10217\,
            I => \N__10208\
        );

    \I__1552\ : Span4Mux_h
    port map (
            O => \N__10214\,
            I => \N__10203\
        );

    \I__1551\ : Span4Mux_h
    port map (
            O => \N__10211\,
            I => \N__10203\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__10208\,
            I => \r_SM_Main_2_N_325_0\
        );

    \I__1549\ : Odrv4
    port map (
            O => \N__10203\,
            I => \r_SM_Main_2_N_325_0\
        );

    \I__1548\ : CascadeMux
    port map (
            O => \N__10198\,
            I => \N__10194\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__10197\,
            I => \N__10190\
        );

    \I__1546\ : InMux
    port map (
            O => \N__10194\,
            I => \N__10187\
        );

    \I__1545\ : InMux
    port map (
            O => \N__10193\,
            I => \N__10184\
        );

    \I__1544\ : InMux
    port map (
            O => \N__10190\,
            I => \N__10181\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__10187\,
            I => \N__10176\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__10184\,
            I => \N__10176\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__10181\,
            I => \N__10173\
        );

    \I__1540\ : Span4Mux_v
    port map (
            O => \N__10176\,
            I => \N__10168\
        );

    \I__1539\ : Span4Mux_h
    port map (
            O => \N__10173\,
            I => \N__10165\
        );

    \I__1538\ : InMux
    port map (
            O => \N__10172\,
            I => \N__10162\
        );

    \I__1537\ : InMux
    port map (
            O => \N__10171\,
            I => \N__10159\
        );

    \I__1536\ : Odrv4
    port map (
            O => \N__10168\,
            I => rx_buf_byte_4
        );

    \I__1535\ : Odrv4
    port map (
            O => \N__10165\,
            I => rx_buf_byte_4
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__10162\,
            I => rx_buf_byte_4
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__10159\,
            I => rx_buf_byte_4
        );

    \I__1532\ : InMux
    port map (
            O => \N__10150\,
            I => \N__10147\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__10147\,
            I => \N__10143\
        );

    \I__1530\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10140\
        );

    \I__1529\ : Span4Mux_h
    port map (
            O => \N__10143\,
            I => \N__10137\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__10140\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_4\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__10137\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_4\
        );

    \I__1526\ : InMux
    port map (
            O => \N__10132\,
            I => \N__10129\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__10129\,
            I => \pc_tx.n6\
        );

    \I__1524\ : ClkMux
    port map (
            O => \N__10126\,
            I => \N__10120\
        );

    \I__1523\ : ClkMux
    port map (
            O => \N__10125\,
            I => \N__10115\
        );

    \I__1522\ : ClkMux
    port map (
            O => \N__10124\,
            I => \N__10108\
        );

    \I__1521\ : ClkMux
    port map (
            O => \N__10123\,
            I => \N__10104\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__10120\,
            I => \N__10101\
        );

    \I__1519\ : ClkMux
    port map (
            O => \N__10119\,
            I => \N__10098\
        );

    \I__1518\ : ClkMux
    port map (
            O => \N__10118\,
            I => \N__10093\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__10115\,
            I => \N__10090\
        );

    \I__1516\ : ClkMux
    port map (
            O => \N__10114\,
            I => \N__10087\
        );

    \I__1515\ : ClkMux
    port map (
            O => \N__10113\,
            I => \N__10084\
        );

    \I__1514\ : ClkMux
    port map (
            O => \N__10112\,
            I => \N__10079\
        );

    \I__1513\ : ClkMux
    port map (
            O => \N__10111\,
            I => \N__10076\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__10108\,
            I => \N__10072\
        );

    \I__1511\ : ClkMux
    port map (
            O => \N__10107\,
            I => \N__10069\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__10104\,
            I => \N__10066\
        );

    \I__1509\ : Span4Mux_v
    port map (
            O => \N__10101\,
            I => \N__10063\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__10098\,
            I => \N__10060\
        );

    \I__1507\ : ClkMux
    port map (
            O => \N__10097\,
            I => \N__10057\
        );

    \I__1506\ : ClkMux
    port map (
            O => \N__10096\,
            I => \N__10054\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__10093\,
            I => \N__10051\
        );

    \I__1504\ : Span4Mux_h
    port map (
            O => \N__10090\,
            I => \N__10048\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__10087\,
            I => \N__10045\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__10084\,
            I => \N__10042\
        );

    \I__1501\ : ClkMux
    port map (
            O => \N__10083\,
            I => \N__10039\
        );

    \I__1500\ : ClkMux
    port map (
            O => \N__10082\,
            I => \N__10036\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__10079\,
            I => \N__10033\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__10076\,
            I => \N__10030\
        );

    \I__1497\ : ClkMux
    port map (
            O => \N__10075\,
            I => \N__10027\
        );

    \I__1496\ : Span4Mux_v
    port map (
            O => \N__10072\,
            I => \N__10020\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__10069\,
            I => \N__10020\
        );

    \I__1494\ : Span4Mux_v
    port map (
            O => \N__10066\,
            I => \N__10017\
        );

    \I__1493\ : Span4Mux_v
    port map (
            O => \N__10063\,
            I => \N__10014\
        );

    \I__1492\ : Span4Mux_h
    port map (
            O => \N__10060\,
            I => \N__10007\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__10057\,
            I => \N__10007\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__10054\,
            I => \N__10007\
        );

    \I__1489\ : Span4Mux_h
    port map (
            O => \N__10051\,
            I => \N__10004\
        );

    \I__1488\ : Span4Mux_h
    port map (
            O => \N__10048\,
            I => \N__9995\
        );

    \I__1487\ : Span4Mux_h
    port map (
            O => \N__10045\,
            I => \N__9995\
        );

    \I__1486\ : Span4Mux_v
    port map (
            O => \N__10042\,
            I => \N__9995\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__10039\,
            I => \N__9995\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__10036\,
            I => \N__9992\
        );

    \I__1483\ : Span4Mux_v
    port map (
            O => \N__10033\,
            I => \N__9985\
        );

    \I__1482\ : Span4Mux_h
    port map (
            O => \N__10030\,
            I => \N__9985\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__10027\,
            I => \N__9985\
        );

    \I__1480\ : InMux
    port map (
            O => \N__10026\,
            I => \N__9982\
        );

    \I__1479\ : ClkMux
    port map (
            O => \N__10025\,
            I => \N__9979\
        );

    \I__1478\ : Span4Mux_v
    port map (
            O => \N__10020\,
            I => \N__9975\
        );

    \I__1477\ : Span4Mux_v
    port map (
            O => \N__10017\,
            I => \N__9968\
        );

    \I__1476\ : Span4Mux_v
    port map (
            O => \N__10014\,
            I => \N__9968\
        );

    \I__1475\ : Span4Mux_v
    port map (
            O => \N__10007\,
            I => \N__9968\
        );

    \I__1474\ : Span4Mux_v
    port map (
            O => \N__10004\,
            I => \N__9961\
        );

    \I__1473\ : Span4Mux_v
    port map (
            O => \N__9995\,
            I => \N__9961\
        );

    \I__1472\ : Span4Mux_h
    port map (
            O => \N__9992\,
            I => \N__9961\
        );

    \I__1471\ : Span4Mux_v
    port map (
            O => \N__9985\,
            I => \N__9956\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__9982\,
            I => \N__9956\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__9979\,
            I => \N__9953\
        );

    \I__1468\ : InMux
    port map (
            O => \N__9978\,
            I => \N__9950\
        );

    \I__1467\ : Odrv4
    port map (
            O => \N__9975\,
            I => \spi0.spi_clk\
        );

    \I__1466\ : Odrv4
    port map (
            O => \N__9968\,
            I => \spi0.spi_clk\
        );

    \I__1465\ : Odrv4
    port map (
            O => \N__9961\,
            I => \spi0.spi_clk\
        );

    \I__1464\ : Odrv4
    port map (
            O => \N__9956\,
            I => \spi0.spi_clk\
        );

    \I__1463\ : Odrv12
    port map (
            O => \N__9953\,
            I => \spi0.spi_clk\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__9950\,
            I => \spi0.spi_clk\
        );

    \I__1461\ : CascadeMux
    port map (
            O => \N__9937\,
            I => \n2446_cascade_\
        );

    \I__1460\ : InMux
    port map (
            O => \N__9934\,
            I => \N__9931\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__9931\,
            I => tx_shift_reg_4
        );

    \I__1458\ : InMux
    port map (
            O => \N__9928\,
            I => \N__9925\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__9925\,
            I => tx_shift_reg_8
        );

    \I__1456\ : InMux
    port map (
            O => \N__9922\,
            I => \N__9919\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__9919\,
            I => tx_shift_reg_3
        );

    \I__1454\ : InMux
    port map (
            O => \N__9916\,
            I => \N__9913\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__9913\,
            I => \N__9910\
        );

    \I__1452\ : Span4Mux_v
    port map (
            O => \N__9910\,
            I => \N__9907\
        );

    \I__1451\ : Sp12to4
    port map (
            O => \N__9907\,
            I => \N__9904\
        );

    \I__1450\ : Odrv12
    port map (
            O => \N__9904\,
            I => \spi0.CS_w\
        );

    \I__1449\ : SRMux
    port map (
            O => \N__9901\,
            I => \N__9898\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__9898\,
            I => \N__9894\
        );

    \I__1447\ : InMux
    port map (
            O => \N__9897\,
            I => \N__9891\
        );

    \I__1446\ : Span4Mux_h
    port map (
            O => \N__9894\,
            I => \N__9888\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__9891\,
            I => \N__9885\
        );

    \I__1444\ : Odrv4
    port map (
            O => \N__9888\,
            I => \spi0.n2715\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__9885\,
            I => \spi0.n2715\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__9880\,
            I => \pc_tx.n5_cascade_\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__9877\,
            I => \pc_tx.n4905_cascade_\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__9874\,
            I => \pc_tx.r_SM_Main_2_N_322_1_cascade_\
        );

    \I__1439\ : InMux
    port map (
            O => \N__9871\,
            I => \N__9867\
        );

    \I__1438\ : InMux
    port map (
            O => \N__9870\,
            I => \N__9864\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__9867\,
            I => \N__9859\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__9864\,
            I => \N__9859\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__9859\,
            I => \pc_tx.n3763\
        );

    \I__1434\ : InMux
    port map (
            O => \N__9856\,
            I => \N__9853\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__9853\,
            I => \pc_tx.n2069\
        );

    \I__1432\ : CEMux
    port map (
            O => \N__9850\,
            I => \N__9847\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__9847\,
            I => \N__9843\
        );

    \I__1430\ : InMux
    port map (
            O => \N__9846\,
            I => \N__9840\
        );

    \I__1429\ : Span4Mux_v
    port map (
            O => \N__9843\,
            I => \N__9834\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__9840\,
            I => \N__9834\
        );

    \I__1427\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9831\
        );

    \I__1426\ : Odrv4
    port map (
            O => \N__9834\,
            I => \pc_tx.n5484\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__9831\,
            I => \pc_tx.n5484\
        );

    \I__1424\ : InMux
    port map (
            O => \N__9826\,
            I => \N__9820\
        );

    \I__1423\ : InMux
    port map (
            O => \N__9825\,
            I => \N__9820\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__9820\,
            I => \spi0.state_next_2__N_453\
        );

    \I__1421\ : InMux
    port map (
            O => \N__9817\,
            I => \N__9812\
        );

    \I__1420\ : InMux
    port map (
            O => \N__9816\,
            I => \N__9809\
        );

    \I__1419\ : InMux
    port map (
            O => \N__9815\,
            I => \N__9806\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__9812\,
            I => \spi0.state_next_2__N_452\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__9809\,
            I => \spi0.state_next_2__N_452\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__9806\,
            I => \spi0.state_next_2__N_452\
        );

    \I__1415\ : CascadeMux
    port map (
            O => \N__9799\,
            I => \spi0.n5561_cascade_\
        );

    \I__1414\ : InMux
    port map (
            O => \N__9796\,
            I => \N__9793\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__9793\,
            I => \spi0.n25\
        );

    \I__1412\ : InMux
    port map (
            O => \N__9790\,
            I => \N__9787\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__9787\,
            I => \spi0.n13\
        );

    \I__1410\ : InMux
    port map (
            O => \N__9784\,
            I => \N__9777\
        );

    \I__1409\ : InMux
    port map (
            O => \N__9783\,
            I => \N__9770\
        );

    \I__1408\ : InMux
    port map (
            O => \N__9782\,
            I => \N__9770\
        );

    \I__1407\ : InMux
    port map (
            O => \N__9781\,
            I => \N__9770\
        );

    \I__1406\ : InMux
    port map (
            O => \N__9780\,
            I => \N__9767\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__9777\,
            I => n982
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__9770\,
            I => n982
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__9767\,
            I => n982
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__9760\,
            I => \N__9756\
        );

    \I__1401\ : InMux
    port map (
            O => \N__9759\,
            I => \N__9752\
        );

    \I__1400\ : InMux
    port map (
            O => \N__9756\,
            I => \N__9747\
        );

    \I__1399\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9747\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__9752\,
            I => \spi0.n2120\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__9747\,
            I => \spi0.n2120\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__9742\,
            I => \spi0.n13_cascade_\
        );

    \I__1395\ : InMux
    port map (
            O => \N__9739\,
            I => \N__9736\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__9736\,
            I => \spi0.state_next_0\
        );

    \I__1393\ : InMux
    port map (
            O => \N__9733\,
            I => \N__9730\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__9730\,
            I => \N__9727\
        );

    \I__1391\ : Odrv4
    port map (
            O => \N__9727\,
            I => \mem_LUT_data_raw_r_5\
        );

    \I__1390\ : InMux
    port map (
            O => \N__9724\,
            I => \N__9721\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__9721\,
            I => \N__9718\
        );

    \I__1388\ : Span4Mux_v
    port map (
            O => \N__9718\,
            I => \N__9714\
        );

    \I__1387\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9711\
        );

    \I__1386\ : Odrv4
    port map (
            O => \N__9714\,
            I => fifo_temp_output_5
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__9711\,
            I => fifo_temp_output_5
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__9706\,
            I => \N__9702\
        );

    \I__1383\ : InMux
    port map (
            O => \N__9705\,
            I => \N__9699\
        );

    \I__1382\ : InMux
    port map (
            O => \N__9702\,
            I => \N__9696\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__9699\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_7\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__9696\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_7\
        );

    \I__1379\ : InMux
    port map (
            O => \N__9691\,
            I => \N__9688\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__9688\,
            I => \N__9685\
        );

    \I__1377\ : Odrv4
    port map (
            O => \N__9685\,
            I => \tx_fifo.lscc_fifo_inst.n5684\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__9682\,
            I => \N__9679\
        );

    \I__1375\ : InMux
    port map (
            O => \N__9679\,
            I => \N__9676\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__9676\,
            I => \N__9673\
        );

    \I__1373\ : Odrv4
    port map (
            O => \N__9673\,
            I => \mem_LUT_data_raw_r_1\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__9670\,
            I => \N__9667\
        );

    \I__1371\ : InMux
    port map (
            O => \N__9667\,
            I => \N__9664\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__9664\,
            I => \N__9660\
        );

    \I__1369\ : InMux
    port map (
            O => \N__9663\,
            I => \N__9657\
        );

    \I__1368\ : Odrv12
    port map (
            O => \N__9660\,
            I => fifo_temp_output_1
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__9657\,
            I => fifo_temp_output_1
        );

    \I__1366\ : InMux
    port map (
            O => \N__9652\,
            I => \N__9649\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__9649\,
            I => \N__9646\
        );

    \I__1364\ : Span4Mux_h
    port map (
            O => \N__9646\,
            I => \N__9643\
        );

    \I__1363\ : Span4Mux_v
    port map (
            O => \N__9643\,
            I => \N__9640\
        );

    \I__1362\ : Span4Mux_v
    port map (
            O => \N__9640\,
            I => \N__9637\
        );

    \I__1361\ : Span4Mux_v
    port map (
            O => \N__9637\,
            I => \N__9634\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__9634\,
            I => \FIFO_D8_c_8\
        );

    \I__1359\ : IoInMux
    port map (
            O => \N__9631\,
            I => \N__9628\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__9628\,
            I => \N__9625\
        );

    \I__1357\ : Span4Mux_s2_h
    port map (
            O => \N__9625\,
            I => \N__9622\
        );

    \I__1356\ : Span4Mux_h
    port map (
            O => \N__9622\,
            I => \N__9619\
        );

    \I__1355\ : Span4Mux_h
    port map (
            O => \N__9619\,
            I => \N__9616\
        );

    \I__1354\ : Sp12to4
    port map (
            O => \N__9616\,
            I => \N__9613\
        );

    \I__1353\ : Span12Mux_v
    port map (
            O => \N__9613\,
            I => \N__9610\
        );

    \I__1352\ : Odrv12
    port map (
            O => \N__9610\,
            I => \DATA8_c_8\
        );

    \I__1351\ : CascadeMux
    port map (
            O => \N__9607\,
            I => \spi0.n5552_cascade_\
        );

    \I__1350\ : CascadeMux
    port map (
            O => \N__9604\,
            I => \spi0.state_next_2_cascade_\
        );

    \I__1349\ : CascadeMux
    port map (
            O => \N__9601\,
            I => \spi0.n4_cascade_\
        );

    \I__1348\ : CascadeMux
    port map (
            O => \N__9598\,
            I => \N__9595\
        );

    \I__1347\ : InMux
    port map (
            O => \N__9595\,
            I => \N__9592\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__9592\,
            I => \spi0.n492\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__9589\,
            I => \N__9586\
        );

    \I__1344\ : InMux
    port map (
            O => \N__9586\,
            I => \N__9583\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__9583\,
            I => \N__9580\
        );

    \I__1342\ : Odrv4
    port map (
            O => \N__9580\,
            I => \spi0.n491\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__9577\,
            I => \N__9572\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__9576\,
            I => \N__9568\
        );

    \I__1339\ : CascadeMux
    port map (
            O => \N__9575\,
            I => \N__9565\
        );

    \I__1338\ : InMux
    port map (
            O => \N__9572\,
            I => \N__9562\
        );

    \I__1337\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9559\
        );

    \I__1336\ : InMux
    port map (
            O => \N__9568\,
            I => \N__9556\
        );

    \I__1335\ : InMux
    port map (
            O => \N__9565\,
            I => \N__9553\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__9562\,
            I => \N__9546\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__9559\,
            I => \N__9546\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__9556\,
            I => \N__9546\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__9553\,
            I => \state_next_2__N_454\
        );

    \I__1330\ : Odrv4
    port map (
            O => \N__9546\,
            I => \state_next_2__N_454\
        );

    \I__1329\ : InMux
    port map (
            O => \N__9541\,
            I => \N__9537\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__9540\,
            I => \N__9534\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__9537\,
            I => \N__9531\
        );

    \I__1326\ : InMux
    port map (
            O => \N__9534\,
            I => \N__9528\
        );

    \I__1325\ : Odrv12
    port map (
            O => \N__9531\,
            I => \spi0.n1005\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__9528\,
            I => \spi0.n1005\
        );

    \I__1323\ : CascadeMux
    port map (
            O => \N__9523\,
            I => \n982_cascade_\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__9520\,
            I => \N__9511\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__9519\,
            I => \N__9508\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__9518\,
            I => \N__9505\
        );

    \I__1319\ : InMux
    port map (
            O => \N__9517\,
            I => \N__9497\
        );

    \I__1318\ : InMux
    port map (
            O => \N__9516\,
            I => \N__9497\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__9515\,
            I => \N__9494\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__9514\,
            I => \N__9487\
        );

    \I__1315\ : InMux
    port map (
            O => \N__9511\,
            I => \N__9473\
        );

    \I__1314\ : InMux
    port map (
            O => \N__9508\,
            I => \N__9473\
        );

    \I__1313\ : InMux
    port map (
            O => \N__9505\,
            I => \N__9473\
        );

    \I__1312\ : InMux
    port map (
            O => \N__9504\,
            I => \N__9473\
        );

    \I__1311\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9473\
        );

    \I__1310\ : InMux
    port map (
            O => \N__9502\,
            I => \N__9473\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__9497\,
            I => \N__9470\
        );

    \I__1308\ : InMux
    port map (
            O => \N__9494\,
            I => \N__9461\
        );

    \I__1307\ : InMux
    port map (
            O => \N__9493\,
            I => \N__9461\
        );

    \I__1306\ : InMux
    port map (
            O => \N__9492\,
            I => \N__9461\
        );

    \I__1305\ : InMux
    port map (
            O => \N__9491\,
            I => \N__9461\
        );

    \I__1304\ : InMux
    port map (
            O => \N__9490\,
            I => \N__9458\
        );

    \I__1303\ : InMux
    port map (
            O => \N__9487\,
            I => \N__9453\
        );

    \I__1302\ : InMux
    port map (
            O => \N__9486\,
            I => \N__9453\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__9473\,
            I => \spi0.state_next_1\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__9470\,
            I => \spi0.state_next_1\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__9461\,
            I => \spi0.state_next_1\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__9458\,
            I => \spi0.state_next_1\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__9453\,
            I => \spi0.state_next_1\
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__9442\,
            I => \N__9439\
        );

    \I__1295\ : InMux
    port map (
            O => \N__9439\,
            I => \N__9436\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__9436\,
            I => \spi0.n495\
        );

    \I__1293\ : InMux
    port map (
            O => \N__9433\,
            I => \N__9426\
        );

    \I__1292\ : InMux
    port map (
            O => \N__9432\,
            I => \N__9407\
        );

    \I__1291\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9407\
        );

    \I__1290\ : InMux
    port map (
            O => \N__9430\,
            I => \N__9407\
        );

    \I__1289\ : InMux
    port map (
            O => \N__9429\,
            I => \N__9407\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__9426\,
            I => \N__9404\
        );

    \I__1287\ : InMux
    port map (
            O => \N__9425\,
            I => \N__9399\
        );

    \I__1286\ : InMux
    port map (
            O => \N__9424\,
            I => \N__9399\
        );

    \I__1285\ : InMux
    port map (
            O => \N__9423\,
            I => \N__9384\
        );

    \I__1284\ : InMux
    port map (
            O => \N__9422\,
            I => \N__9384\
        );

    \I__1283\ : InMux
    port map (
            O => \N__9421\,
            I => \N__9384\
        );

    \I__1282\ : InMux
    port map (
            O => \N__9420\,
            I => \N__9384\
        );

    \I__1281\ : InMux
    port map (
            O => \N__9419\,
            I => \N__9384\
        );

    \I__1280\ : InMux
    port map (
            O => \N__9418\,
            I => \N__9384\
        );

    \I__1279\ : InMux
    port map (
            O => \N__9417\,
            I => \N__9384\
        );

    \I__1278\ : InMux
    port map (
            O => \N__9416\,
            I => \N__9381\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__9407\,
            I => \spi0.n4\
        );

    \I__1276\ : Odrv4
    port map (
            O => \N__9404\,
            I => \spi0.n4\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__9399\,
            I => \spi0.n4\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__9384\,
            I => \spi0.n4\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__9381\,
            I => \spi0.n4\
        );

    \I__1272\ : InMux
    port map (
            O => \N__9370\,
            I => \N__9367\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__9367\,
            I => \N__9364\
        );

    \I__1270\ : Span4Mux_h
    port map (
            O => \N__9364\,
            I => \N__9361\
        );

    \I__1269\ : Odrv4
    port map (
            O => \N__9361\,
            I => \mem_LUT_data_raw_r_3\
        );

    \I__1268\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9355\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__9355\,
            I => \N__9351\
        );

    \I__1266\ : InMux
    port map (
            O => \N__9354\,
            I => \N__9348\
        );

    \I__1265\ : Odrv4
    port map (
            O => \N__9351\,
            I => fifo_temp_output_3
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__9348\,
            I => fifo_temp_output_3
        );

    \I__1263\ : CascadeMux
    port map (
            O => \N__9343\,
            I => \N__9340\
        );

    \I__1262\ : InMux
    port map (
            O => \N__9340\,
            I => \N__9337\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__9337\,
            I => \N__9334\
        );

    \I__1260\ : Span4Mux_h
    port map (
            O => \N__9334\,
            I => \N__9331\
        );

    \I__1259\ : Odrv4
    port map (
            O => \N__9331\,
            I => \mem_LUT_data_raw_r_0\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__9328\,
            I => \N__9324\
        );

    \I__1257\ : InMux
    port map (
            O => \N__9327\,
            I => \N__9317\
        );

    \I__1256\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9317\
        );

    \I__1255\ : InMux
    port map (
            O => \N__9323\,
            I => \N__9314\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__9322\,
            I => \N__9311\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__9317\,
            I => \N__9308\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__9314\,
            I => \N__9305\
        );

    \I__1251\ : InMux
    port map (
            O => \N__9311\,
            I => \N__9302\
        );

    \I__1250\ : Span4Mux_v
    port map (
            O => \N__9308\,
            I => \N__9298\
        );

    \I__1249\ : Span4Mux_h
    port map (
            O => \N__9305\,
            I => \N__9295\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__9302\,
            I => \N__9292\
        );

    \I__1247\ : InMux
    port map (
            O => \N__9301\,
            I => \N__9289\
        );

    \I__1246\ : Odrv4
    port map (
            O => \N__9298\,
            I => rx_buf_byte_1
        );

    \I__1245\ : Odrv4
    port map (
            O => \N__9295\,
            I => rx_buf_byte_1
        );

    \I__1244\ : Odrv12
    port map (
            O => \N__9292\,
            I => rx_buf_byte_1
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__9289\,
            I => rx_buf_byte_1
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__9280\,
            I => \N__9276\
        );

    \I__1241\ : InMux
    port map (
            O => \N__9279\,
            I => \N__9273\
        );

    \I__1240\ : InMux
    port map (
            O => \N__9276\,
            I => \N__9270\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__9273\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_1\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__9270\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_1\
        );

    \I__1237\ : InMux
    port map (
            O => \N__9265\,
            I => \N__9259\
        );

    \I__1236\ : InMux
    port map (
            O => \N__9264\,
            I => \N__9259\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__9259\,
            I => \r_Tx_Data_1\
        );

    \I__1234\ : InMux
    port map (
            O => \N__9256\,
            I => \N__9252\
        );

    \I__1233\ : InMux
    port map (
            O => \N__9255\,
            I => \N__9249\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__9252\,
            I => \N__9246\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__9249\,
            I => fifo_temp_output_0
        );

    \I__1230\ : Odrv4
    port map (
            O => \N__9246\,
            I => fifo_temp_output_0
        );

    \I__1229\ : InMux
    port map (
            O => \N__9241\,
            I => \N__9232\
        );

    \I__1228\ : InMux
    port map (
            O => \N__9240\,
            I => \N__9227\
        );

    \I__1227\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9227\
        );

    \I__1226\ : InMux
    port map (
            O => \N__9238\,
            I => \N__9222\
        );

    \I__1225\ : InMux
    port map (
            O => \N__9237\,
            I => \N__9222\
        );

    \I__1224\ : InMux
    port map (
            O => \N__9236\,
            I => \N__9217\
        );

    \I__1223\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9217\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__9232\,
            I => n2366
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__9227\,
            I => n2366
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__9222\,
            I => n2366
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__9217\,
            I => n2366
        );

    \I__1218\ : InMux
    port map (
            O => \N__9208\,
            I => \N__9202\
        );

    \I__1217\ : InMux
    port map (
            O => \N__9207\,
            I => \N__9202\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__9202\,
            I => \r_Tx_Data_0\
        );

    \I__1215\ : InMux
    port map (
            O => \N__9199\,
            I => \N__9195\
        );

    \I__1214\ : InMux
    port map (
            O => \N__9198\,
            I => \N__9192\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__9195\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_4\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__9192\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_4\
        );

    \I__1211\ : CascadeMux
    port map (
            O => \N__9187\,
            I => \spi0.n2120_cascade_\
        );

    \I__1210\ : InMux
    port map (
            O => \N__9184\,
            I => \N__9181\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__9181\,
            I => \spi0.n5552\
        );

    \I__1208\ : InMux
    port map (
            O => \N__9178\,
            I => \N__9174\
        );

    \I__1207\ : InMux
    port map (
            O => \N__9177\,
            I => \N__9171\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__9174\,
            I => \r_Tx_Data_6\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__9171\,
            I => \r_Tx_Data_6\
        );

    \I__1204\ : InMux
    port map (
            O => \N__9166\,
            I => \N__9158\
        );

    \I__1203\ : InMux
    port map (
            O => \N__9165\,
            I => \N__9158\
        );

    \I__1202\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9155\
        );

    \I__1201\ : InMux
    port map (
            O => \N__9163\,
            I => \N__9152\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__9158\,
            I => \pc_tx.r_Bit_Index_1\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__9155\,
            I => \pc_tx.r_Bit_Index_1\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__9152\,
            I => \pc_tx.r_Bit_Index_1\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__9145\,
            I => \pc_tx.n5512_cascade_\
        );

    \I__1196\ : InMux
    port map (
            O => \N__9142\,
            I => \N__9139\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__9139\,
            I => \pc_tx.n5511\
        );

    \I__1194\ : InMux
    port map (
            O => \N__9136\,
            I => \N__9130\
        );

    \I__1193\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9127\
        );

    \I__1192\ : InMux
    port map (
            O => \N__9134\,
            I => \N__9124\
        );

    \I__1191\ : InMux
    port map (
            O => \N__9133\,
            I => \N__9121\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__9130\,
            I => \pc_tx.r_Bit_Index_2\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__9127\,
            I => \pc_tx.r_Bit_Index_2\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__9124\,
            I => \pc_tx.r_Bit_Index_2\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__9121\,
            I => \pc_tx.r_Bit_Index_2\
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__9112\,
            I => \pc_tx.n5654_cascade_\
        );

    \I__1185\ : InMux
    port map (
            O => \N__9109\,
            I => \N__9106\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__9106\,
            I => \pc_tx.n5509\
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__9103\,
            I => \pc_tx.o_Tx_Serial_N_354_cascade_\
        );

    \I__1182\ : IoInMux
    port map (
            O => \N__9100\,
            I => \N__9097\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__9097\,
            I => \N__9094\
        );

    \I__1180\ : Span12Mux_s7_h
    port map (
            O => \N__9094\,
            I => \N__9091\
        );

    \I__1179\ : Span12Mux_h
    port map (
            O => \N__9091\,
            I => \N__9088\
        );

    \I__1178\ : Odrv12
    port map (
            O => \N__9088\,
            I => \pc_tx.n3_adj_632\
        );

    \I__1177\ : SRMux
    port map (
            O => \N__9085\,
            I => \N__9082\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__9082\,
            I => \pc_tx.n5486\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__9079\,
            I => \n2366_cascade_\
        );

    \I__1174\ : InMux
    port map (
            O => \N__9076\,
            I => \N__9070\
        );

    \I__1173\ : InMux
    port map (
            O => \N__9075\,
            I => \N__9070\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__9070\,
            I => \r_Tx_Data_7\
        );

    \I__1171\ : InMux
    port map (
            O => \N__9067\,
            I => \N__9055\
        );

    \I__1170\ : InMux
    port map (
            O => \N__9066\,
            I => \N__9055\
        );

    \I__1169\ : InMux
    port map (
            O => \N__9065\,
            I => \N__9050\
        );

    \I__1168\ : InMux
    port map (
            O => \N__9064\,
            I => \N__9050\
        );

    \I__1167\ : InMux
    port map (
            O => \N__9063\,
            I => \N__9047\
        );

    \I__1166\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9044\
        );

    \I__1165\ : InMux
    port map (
            O => \N__9061\,
            I => \N__9039\
        );

    \I__1164\ : InMux
    port map (
            O => \N__9060\,
            I => \N__9039\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__9055\,
            I => \pc_tx.r_Bit_Index_0\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__9050\,
            I => \pc_tx.r_Bit_Index_0\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__9047\,
            I => \pc_tx.r_Bit_Index_0\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__9044\,
            I => \pc_tx.r_Bit_Index_0\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__9039\,
            I => \pc_tx.r_Bit_Index_0\
        );

    \I__1158\ : InMux
    port map (
            O => \N__9028\,
            I => \N__9025\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__9025\,
            I => \pc_tx.n5508\
        );

    \I__1156\ : InMux
    port map (
            O => \N__9022\,
            I => \N__9018\
        );

    \I__1155\ : InMux
    port map (
            O => \N__9021\,
            I => \N__9015\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__9018\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_4\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__9015\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_4\
        );

    \I__1152\ : CascadeMux
    port map (
            O => \N__9010\,
            I => \N__9007\
        );

    \I__1151\ : InMux
    port map (
            O => \N__9007\,
            I => \N__9004\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__9004\,
            I => \N__9001\
        );

    \I__1149\ : Odrv4
    port map (
            O => \N__9001\,
            I => \mem_LUT_data_raw_r_2\
        );

    \I__1148\ : InMux
    port map (
            O => \N__8998\,
            I => \N__8994\
        );

    \I__1147\ : InMux
    port map (
            O => \N__8997\,
            I => \N__8991\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__8994\,
            I => fifo_temp_output_4
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__8991\,
            I => fifo_temp_output_4
        );

    \I__1144\ : InMux
    port map (
            O => \N__8986\,
            I => \N__8982\
        );

    \I__1143\ : InMux
    port map (
            O => \N__8985\,
            I => \N__8979\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__8982\,
            I => fifo_temp_output_2
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__8979\,
            I => fifo_temp_output_2
        );

    \I__1140\ : InMux
    port map (
            O => \N__8974\,
            I => \N__8968\
        );

    \I__1139\ : InMux
    port map (
            O => \N__8973\,
            I => \N__8968\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__8968\,
            I => \r_Tx_Data_3\
        );

    \I__1137\ : InMux
    port map (
            O => \N__8965\,
            I => \N__8959\
        );

    \I__1136\ : InMux
    port map (
            O => \N__8964\,
            I => \N__8959\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__8959\,
            I => \r_Tx_Data_2\
        );

    \I__1134\ : InMux
    port map (
            O => \N__8956\,
            I => \N__8950\
        );

    \I__1133\ : InMux
    port map (
            O => \N__8955\,
            I => \N__8950\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__8950\,
            I => \r_Tx_Data_5\
        );

    \I__1131\ : InMux
    port map (
            O => \N__8947\,
            I => \N__8941\
        );

    \I__1130\ : InMux
    port map (
            O => \N__8946\,
            I => \N__8941\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__8941\,
            I => \r_Tx_Data_4\
        );

    \I__1128\ : InMux
    port map (
            O => \N__8938\,
            I => \N__8935\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__8935\,
            I => n5414
        );

    \I__1126\ : InMux
    port map (
            O => \N__8932\,
            I => \N__8928\
        );

    \I__1125\ : InMux
    port map (
            O => \N__8931\,
            I => \N__8925\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__8928\,
            I => \spi0.spi_clk_counter_0\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__8925\,
            I => \spi0.spi_clk_counter_0\
        );

    \I__1122\ : InMux
    port map (
            O => \N__8920\,
            I => \bfn_8_12_0_\
        );

    \I__1121\ : InMux
    port map (
            O => \N__8917\,
            I => \N__8913\
        );

    \I__1120\ : InMux
    port map (
            O => \N__8916\,
            I => \N__8910\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__8913\,
            I => \spi0.spi_clk_counter_1\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__8910\,
            I => \spi0.spi_clk_counter_1\
        );

    \I__1117\ : InMux
    port map (
            O => \N__8905\,
            I => \spi0.n4874\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__8902\,
            I => \N__8899\
        );

    \I__1115\ : InMux
    port map (
            O => \N__8899\,
            I => \N__8895\
        );

    \I__1114\ : InMux
    port map (
            O => \N__8898\,
            I => \N__8892\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__8895\,
            I => \spi0.spi_clk_counter_2\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__8892\,
            I => \spi0.spi_clk_counter_2\
        );

    \I__1111\ : InMux
    port map (
            O => \N__8887\,
            I => \spi0.n4875\
        );

    \I__1110\ : InMux
    port map (
            O => \N__8884\,
            I => \N__8880\
        );

    \I__1109\ : InMux
    port map (
            O => \N__8883\,
            I => \N__8877\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__8880\,
            I => \spi0.spi_clk_counter_3\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__8877\,
            I => \spi0.spi_clk_counter_3\
        );

    \I__1106\ : InMux
    port map (
            O => \N__8872\,
            I => \spi0.n4876\
        );

    \I__1105\ : CascadeMux
    port map (
            O => \N__8869\,
            I => \N__8866\
        );

    \I__1104\ : InMux
    port map (
            O => \N__8866\,
            I => \N__8862\
        );

    \I__1103\ : InMux
    port map (
            O => \N__8865\,
            I => \N__8859\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__8862\,
            I => \spi0.spi_clk_counter_4\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__8859\,
            I => \spi0.spi_clk_counter_4\
        );

    \I__1100\ : InMux
    port map (
            O => \N__8854\,
            I => \spi0.n4877\
        );

    \I__1099\ : InMux
    port map (
            O => \N__8851\,
            I => \N__8847\
        );

    \I__1098\ : InMux
    port map (
            O => \N__8850\,
            I => \N__8844\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__8847\,
            I => \spi0.spi_clk_counter_5\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__8844\,
            I => \spi0.spi_clk_counter_5\
        );

    \I__1095\ : InMux
    port map (
            O => \N__8839\,
            I => \spi0.n4878\
        );

    \I__1094\ : CascadeMux
    port map (
            O => \N__8836\,
            I => \N__8833\
        );

    \I__1093\ : InMux
    port map (
            O => \N__8833\,
            I => \N__8829\
        );

    \I__1092\ : InMux
    port map (
            O => \N__8832\,
            I => \N__8826\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__8829\,
            I => \spi0.spi_clk_counter_6\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__8826\,
            I => \spi0.spi_clk_counter_6\
        );

    \I__1089\ : InMux
    port map (
            O => \N__8821\,
            I => \spi0.n4879\
        );

    \I__1088\ : InMux
    port map (
            O => \N__8818\,
            I => \spi0.n4880\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__8815\,
            I => \N__8811\
        );

    \I__1086\ : InMux
    port map (
            O => \N__8814\,
            I => \N__8808\
        );

    \I__1085\ : InMux
    port map (
            O => \N__8811\,
            I => \N__8805\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__8808\,
            I => \spi0.spi_clk_counter_7\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__8805\,
            I => \spi0.spi_clk_counter_7\
        );

    \I__1082\ : InMux
    port map (
            O => \N__8800\,
            I => \N__8797\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__8797\,
            I => \N__8794\
        );

    \I__1080\ : Span12Mux_v
    port map (
            O => \N__8794\,
            I => \N__8791\
        );

    \I__1079\ : Span12Mux_v
    port map (
            O => \N__8791\,
            I => \N__8788\
        );

    \I__1078\ : Odrv12
    port map (
            O => \N__8788\,
            I => \FIFO_D18_c_18\
        );

    \I__1077\ : IoInMux
    port map (
            O => \N__8785\,
            I => \N__8782\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__8782\,
            I => \N__8779\
        );

    \I__1075\ : Span12Mux_s11_v
    port map (
            O => \N__8779\,
            I => \N__8776\
        );

    \I__1074\ : Span12Mux_h
    port map (
            O => \N__8776\,
            I => \N__8773\
        );

    \I__1073\ : Odrv12
    port map (
            O => \N__8773\,
            I => \DATA18_c_18\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__8770\,
            I => \N__8766\
        );

    \I__1071\ : InMux
    port map (
            O => \N__8769\,
            I => \N__8763\
        );

    \I__1070\ : InMux
    port map (
            O => \N__8766\,
            I => \N__8760\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__8763\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_7\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__8760\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_7\
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__8755\,
            I => \N__8751\
        );

    \I__1066\ : InMux
    port map (
            O => \N__8754\,
            I => \N__8748\
        );

    \I__1065\ : InMux
    port map (
            O => \N__8751\,
            I => \N__8745\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__8748\,
            I => \N__8742\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__8745\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_7\
        );

    \I__1062\ : Odrv4
    port map (
            O => \N__8742\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_7\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__8737\,
            I => \N__8733\
        );

    \I__1060\ : InMux
    port map (
            O => \N__8736\,
            I => \N__8730\
        );

    \I__1059\ : InMux
    port map (
            O => \N__8733\,
            I => \N__8727\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__8730\,
            I => \N__8724\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__8727\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_4\
        );

    \I__1056\ : Odrv12
    port map (
            O => \N__8724\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_4\
        );

    \I__1055\ : CascadeMux
    port map (
            O => \N__8719\,
            I => \spi0.n14_cascade_\
        );

    \I__1054\ : InMux
    port map (
            O => \N__8716\,
            I => \N__8713\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__8713\,
            I => \N__8709\
        );

    \I__1052\ : InMux
    port map (
            O => \N__8712\,
            I => \N__8706\
        );

    \I__1051\ : Odrv4
    port map (
            O => \N__8709\,
            I => rx_shift_reg_5
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__8706\,
            I => rx_shift_reg_5
        );

    \I__1049\ : InMux
    port map (
            O => \N__8701\,
            I => \N__8694\
        );

    \I__1048\ : InMux
    port map (
            O => \N__8700\,
            I => \N__8694\
        );

    \I__1047\ : InMux
    port map (
            O => \N__8699\,
            I => \N__8691\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__8694\,
            I => \N__8688\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__8691\,
            I => \N__8685\
        );

    \I__1044\ : Span12Mux_v
    port map (
            O => \N__8688\,
            I => \N__8677\
        );

    \I__1043\ : Span4Mux_h
    port map (
            O => \N__8685\,
            I => \N__8674\
        );

    \I__1042\ : InMux
    port map (
            O => \N__8684\,
            I => \N__8665\
        );

    \I__1041\ : InMux
    port map (
            O => \N__8683\,
            I => \N__8665\
        );

    \I__1040\ : InMux
    port map (
            O => \N__8682\,
            I => \N__8665\
        );

    \I__1039\ : InMux
    port map (
            O => \N__8681\,
            I => \N__8665\
        );

    \I__1038\ : InMux
    port map (
            O => \N__8680\,
            I => \N__8662\
        );

    \I__1037\ : Odrv12
    port map (
            O => \N__8677\,
            I => \rx_shift_reg_15__N_461\
        );

    \I__1036\ : Odrv4
    port map (
            O => \N__8674\,
            I => \rx_shift_reg_15__N_461\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__8665\,
            I => \rx_shift_reg_15__N_461\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__8662\,
            I => \rx_shift_reg_15__N_461\
        );

    \I__1033\ : InMux
    port map (
            O => \N__8653\,
            I => \N__8650\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__8650\,
            I => \spi0.n10\
        );

    \I__1031\ : InMux
    port map (
            O => \N__8647\,
            I => \N__8644\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__8644\,
            I => \spi0.n483\
        );

    \I__1029\ : CascadeMux
    port map (
            O => \N__8641\,
            I => \N__8638\
        );

    \I__1028\ : InMux
    port map (
            O => \N__8638\,
            I => \N__8635\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__8635\,
            I => \spi0.n484\
        );

    \I__1026\ : InMux
    port map (
            O => \N__8632\,
            I => \N__8629\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__8629\,
            I => \spi0.n485\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__8626\,
            I => \N__8623\
        );

    \I__1023\ : InMux
    port map (
            O => \N__8623\,
            I => \N__8620\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__8620\,
            I => \spi0.n490\
        );

    \I__1021\ : InMux
    port map (
            O => \N__8617\,
            I => \N__8614\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__8614\,
            I => \spi0.n488\
        );

    \I__1019\ : CascadeMux
    port map (
            O => \N__8611\,
            I => \N__8608\
        );

    \I__1018\ : InMux
    port map (
            O => \N__8608\,
            I => \N__8605\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__8605\,
            I => \spi0.n487\
        );

    \I__1016\ : CascadeMux
    port map (
            O => \N__8602\,
            I => \N__8599\
        );

    \I__1015\ : InMux
    port map (
            O => \N__8599\,
            I => \N__8596\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__8596\,
            I => \spi0.n486\
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__8593\,
            I => \N__8590\
        );

    \I__1012\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8587\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__8587\,
            I => \N__8583\
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__8586\,
            I => \N__8578\
        );

    \I__1009\ : Span4Mux_v
    port map (
            O => \N__8583\,
            I => \N__8574\
        );

    \I__1008\ : InMux
    port map (
            O => \N__8582\,
            I => \N__8571\
        );

    \I__1007\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8568\
        );

    \I__1006\ : InMux
    port map (
            O => \N__8578\,
            I => \N__8565\
        );

    \I__1005\ : InMux
    port map (
            O => \N__8577\,
            I => \N__8562\
        );

    \I__1004\ : Odrv4
    port map (
            O => \N__8574\,
            I => rx_buf_byte_6
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__8571\,
            I => rx_buf_byte_6
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__8568\,
            I => rx_buf_byte_6
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__8565\,
            I => rx_buf_byte_6
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__8562\,
            I => rx_buf_byte_6
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__8551\,
            I => \N__8547\
        );

    \I__998\ : InMux
    port map (
            O => \N__8550\,
            I => \N__8544\
        );

    \I__997\ : InMux
    port map (
            O => \N__8547\,
            I => \N__8541\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__8544\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_6\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__8541\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_6\
        );

    \I__994\ : InMux
    port map (
            O => \N__8536\,
            I => \N__8532\
        );

    \I__993\ : InMux
    port map (
            O => \N__8535\,
            I => \N__8529\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__8532\,
            I => \N__8526\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__8529\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_1\
        );

    \I__990\ : Odrv4
    port map (
            O => \N__8526\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_1\
        );

    \I__989\ : CascadeMux
    port map (
            O => \N__8521\,
            I => \N__8518\
        );

    \I__988\ : InMux
    port map (
            O => \N__8518\,
            I => \N__8515\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__8515\,
            I => \N__8511\
        );

    \I__986\ : InMux
    port map (
            O => \N__8514\,
            I => \N__8508\
        );

    \I__985\ : Span4Mux_h
    port map (
            O => \N__8511\,
            I => \N__8505\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__8508\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_1\
        );

    \I__983\ : Odrv4
    port map (
            O => \N__8505\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_1\
        );

    \I__982\ : InMux
    port map (
            O => \N__8500\,
            I => \N__8496\
        );

    \I__981\ : InMux
    port map (
            O => \N__8499\,
            I => \N__8493\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__8496\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_1\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__8493\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_1\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__8488\,
            I => \tx_fifo.lscc_fifo_inst.n5672_cascade_\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__8485\,
            I => \tx_fifo.lscc_fifo_inst.n5678_cascade_\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__8482\,
            I => \N__8479\
        );

    \I__975\ : InMux
    port map (
            O => \N__8479\,
            I => \N__8476\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__8476\,
            I => \mem_LUT_data_raw_r_4\
        );

    \I__973\ : InMux
    port map (
            O => \N__8473\,
            I => \N__8470\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__8470\,
            I => \spi0.n480\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__8467\,
            I => \spi0.state_next_1_cascade_\
        );

    \I__970\ : InMux
    port map (
            O => \N__8464\,
            I => \N__8461\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__8461\,
            I => \spi0.n481\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__8458\,
            I => \N__8455\
        );

    \I__967\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8452\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__8452\,
            I => \spi0.n482\
        );

    \I__965\ : InMux
    port map (
            O => \N__8449\,
            I => \N__8446\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__8446\,
            I => \N__8440\
        );

    \I__963\ : InMux
    port map (
            O => \N__8445\,
            I => \N__8435\
        );

    \I__962\ : InMux
    port map (
            O => \N__8444\,
            I => \N__8435\
        );

    \I__961\ : InMux
    port map (
            O => \N__8443\,
            I => \N__8432\
        );

    \I__960\ : Span4Mux_v
    port map (
            O => \N__8440\,
            I => \N__8428\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__8435\,
            I => \N__8423\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__8432\,
            I => \N__8423\
        );

    \I__957\ : InMux
    port map (
            O => \N__8431\,
            I => \N__8420\
        );

    \I__956\ : Odrv4
    port map (
            O => \N__8428\,
            I => rx_buf_byte_2
        );

    \I__955\ : Odrv12
    port map (
            O => \N__8423\,
            I => rx_buf_byte_2
        );

    \I__954\ : LocalMux
    port map (
            O => \N__8420\,
            I => rx_buf_byte_2
        );

    \I__953\ : CascadeMux
    port map (
            O => \N__8413\,
            I => \N__8409\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__8412\,
            I => \N__8406\
        );

    \I__951\ : InMux
    port map (
            O => \N__8409\,
            I => \N__8403\
        );

    \I__950\ : InMux
    port map (
            O => \N__8406\,
            I => \N__8400\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__8403\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_2\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__8400\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_2\
        );

    \I__947\ : InMux
    port map (
            O => \N__8395\,
            I => \N__8392\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__8392\,
            I => \N__8389\
        );

    \I__945\ : Span4Mux_h
    port map (
            O => \N__8389\,
            I => \N__8385\
        );

    \I__944\ : InMux
    port map (
            O => \N__8388\,
            I => \N__8382\
        );

    \I__943\ : Odrv4
    port map (
            O => \N__8385\,
            I => fifo_temp_output_6
        );

    \I__942\ : LocalMux
    port map (
            O => \N__8382\,
            I => fifo_temp_output_6
        );

    \I__941\ : CascadeMux
    port map (
            O => \N__8377\,
            I => \pc_tx.n3763_cascade_\
        );

    \I__940\ : InMux
    port map (
            O => \N__8374\,
            I => \N__8370\
        );

    \I__939\ : CascadeMux
    port map (
            O => \N__8373\,
            I => \N__8367\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__8370\,
            I => \N__8364\
        );

    \I__937\ : InMux
    port map (
            O => \N__8367\,
            I => \N__8361\
        );

    \I__936\ : Span4Mux_h
    port map (
            O => \N__8364\,
            I => \N__8358\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__8361\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_2\
        );

    \I__934\ : Odrv4
    port map (
            O => \N__8358\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_2\
        );

    \I__933\ : InMux
    port map (
            O => \N__8353\,
            I => \N__8350\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__8350\,
            I => \tx_fifo.lscc_fifo_inst.n5660\
        );

    \I__931\ : InMux
    port map (
            O => \N__8347\,
            I => \N__8343\
        );

    \I__930\ : InMux
    port map (
            O => \N__8346\,
            I => \N__8340\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__8343\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_2\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__8340\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_2\
        );

    \I__927\ : InMux
    port map (
            O => \N__8335\,
            I => \N__8329\
        );

    \I__926\ : InMux
    port map (
            O => \N__8334\,
            I => \N__8329\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__8329\,
            I => \N__8323\
        );

    \I__924\ : InMux
    port map (
            O => \N__8328\,
            I => \N__8320\
        );

    \I__923\ : InMux
    port map (
            O => \N__8327\,
            I => \N__8317\
        );

    \I__922\ : InMux
    port map (
            O => \N__8326\,
            I => \N__8314\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__8323\,
            I => rx_buf_byte_5
        );

    \I__920\ : LocalMux
    port map (
            O => \N__8320\,
            I => rx_buf_byte_5
        );

    \I__919\ : LocalMux
    port map (
            O => \N__8317\,
            I => rx_buf_byte_5
        );

    \I__918\ : LocalMux
    port map (
            O => \N__8314\,
            I => rx_buf_byte_5
        );

    \I__917\ : InMux
    port map (
            O => \N__8305\,
            I => \N__8302\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__8302\,
            I => \N__8298\
        );

    \I__915\ : InMux
    port map (
            O => \N__8301\,
            I => \N__8295\
        );

    \I__914\ : Odrv4
    port map (
            O => \N__8298\,
            I => rx_shift_reg_4
        );

    \I__913\ : LocalMux
    port map (
            O => \N__8295\,
            I => rx_shift_reg_4
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__8290\,
            I => \N__8286\
        );

    \I__911\ : CascadeMux
    port map (
            O => \N__8289\,
            I => \N__8282\
        );

    \I__910\ : InMux
    port map (
            O => \N__8286\,
            I => \N__8276\
        );

    \I__909\ : InMux
    port map (
            O => \N__8285\,
            I => \N__8276\
        );

    \I__908\ : InMux
    port map (
            O => \N__8282\,
            I => \N__8271\
        );

    \I__907\ : InMux
    port map (
            O => \N__8281\,
            I => \N__8271\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__8276\,
            I => \N__8265\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__8271\,
            I => \N__8265\
        );

    \I__904\ : InMux
    port map (
            O => \N__8270\,
            I => \N__8262\
        );

    \I__903\ : Odrv4
    port map (
            O => \N__8265\,
            I => rx_buf_byte_3
        );

    \I__902\ : LocalMux
    port map (
            O => \N__8262\,
            I => rx_buf_byte_3
        );

    \I__901\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8254\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__8254\,
            I => \N__8250\
        );

    \I__899\ : InMux
    port map (
            O => \N__8253\,
            I => \N__8247\
        );

    \I__898\ : Odrv12
    port map (
            O => \N__8250\,
            I => rx_shift_reg_1
        );

    \I__897\ : LocalMux
    port map (
            O => \N__8247\,
            I => rx_shift_reg_1
        );

    \I__896\ : InMux
    port map (
            O => \N__8242\,
            I => \N__8236\
        );

    \I__895\ : InMux
    port map (
            O => \N__8241\,
            I => \N__8236\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__8236\,
            I => rx_shift_reg_2
        );

    \I__893\ : InMux
    port map (
            O => \N__8233\,
            I => \N__8229\
        );

    \I__892\ : InMux
    port map (
            O => \N__8232\,
            I => \N__8226\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__8229\,
            I => rx_shift_reg_3
        );

    \I__890\ : LocalMux
    port map (
            O => \N__8226\,
            I => rx_shift_reg_3
        );

    \I__889\ : IoInMux
    port map (
            O => \N__8221\,
            I => \N__8218\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__8218\,
            I => \N__8215\
        );

    \I__887\ : IoSpan4Mux
    port map (
            O => \N__8215\,
            I => \N__8212\
        );

    \I__886\ : Span4Mux_s1_v
    port map (
            O => \N__8212\,
            I => \N__8209\
        );

    \I__885\ : Sp12to4
    port map (
            O => \N__8209\,
            I => \N__8206\
        );

    \I__884\ : Span12Mux_v
    port map (
            O => \N__8206\,
            I => \N__8202\
        );

    \I__883\ : InMux
    port map (
            O => \N__8205\,
            I => \N__8199\
        );

    \I__882\ : Odrv12
    port map (
            O => \N__8202\,
            I => \SEN_c\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__8199\,
            I => \SEN_c\
        );

    \I__880\ : InMux
    port map (
            O => \N__8194\,
            I => \N__8191\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__8191\,
            I => \N__8188\
        );

    \I__878\ : Span4Mux_v
    port map (
            O => \N__8188\,
            I => \N__8185\
        );

    \I__877\ : Sp12to4
    port map (
            O => \N__8185\,
            I => \N__8182\
        );

    \I__876\ : Span12Mux_h
    port map (
            O => \N__8182\,
            I => \N__8179\
        );

    \I__875\ : Span12Mux_v
    port map (
            O => \N__8179\,
            I => \N__8176\
        );

    \I__874\ : Odrv12
    port map (
            O => \N__8176\,
            I => \FIFO_D25_c_25\
        );

    \I__873\ : IoInMux
    port map (
            O => \N__8173\,
            I => \N__8170\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__8170\,
            I => \N__8167\
        );

    \I__871\ : Span4Mux_s3_v
    port map (
            O => \N__8167\,
            I => \N__8164\
        );

    \I__870\ : Span4Mux_v
    port map (
            O => \N__8164\,
            I => \N__8161\
        );

    \I__869\ : Span4Mux_v
    port map (
            O => \N__8161\,
            I => \N__8158\
        );

    \I__868\ : Sp12to4
    port map (
            O => \N__8158\,
            I => \N__8155\
        );

    \I__867\ : Odrv12
    port map (
            O => \N__8155\,
            I => \DATA25_c_25\
        );

    \I__866\ : InMux
    port map (
            O => \N__8152\,
            I => \N__8149\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__8149\,
            I => \N__8146\
        );

    \I__864\ : Span4Mux_v
    port map (
            O => \N__8146\,
            I => \N__8143\
        );

    \I__863\ : Sp12to4
    port map (
            O => \N__8143\,
            I => \N__8140\
        );

    \I__862\ : Odrv12
    port map (
            O => \N__8140\,
            I => \FIFO_D29_c_29\
        );

    \I__861\ : IoInMux
    port map (
            O => \N__8137\,
            I => \N__8134\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__8134\,
            I => \N__8131\
        );

    \I__859\ : Span4Mux_s3_v
    port map (
            O => \N__8131\,
            I => \N__8128\
        );

    \I__858\ : Span4Mux_v
    port map (
            O => \N__8128\,
            I => \N__8125\
        );

    \I__857\ : Span4Mux_v
    port map (
            O => \N__8125\,
            I => \N__8122\
        );

    \I__856\ : Odrv4
    port map (
            O => \N__8122\,
            I => \DATA29_c_29\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__8119\,
            I => \N__8115\
        );

    \I__854\ : InMux
    port map (
            O => \N__8118\,
            I => \N__8112\
        );

    \I__853\ : InMux
    port map (
            O => \N__8115\,
            I => \N__8109\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__8112\,
            I => \N__8106\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__8109\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_5\
        );

    \I__850\ : Odrv4
    port map (
            O => \N__8106\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_5\
        );

    \I__849\ : CascadeMux
    port map (
            O => \N__8101\,
            I => \N__8097\
        );

    \I__848\ : InMux
    port map (
            O => \N__8100\,
            I => \N__8094\
        );

    \I__847\ : InMux
    port map (
            O => \N__8097\,
            I => \N__8091\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__8094\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_5\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__8091\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_5\
        );

    \I__844\ : InMux
    port map (
            O => \N__8086\,
            I => \N__8082\
        );

    \I__843\ : InMux
    port map (
            O => \N__8085\,
            I => \N__8079\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__8082\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_3\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__8079\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_3\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__8074\,
            I => \N__8070\
        );

    \I__839\ : InMux
    port map (
            O => \N__8073\,
            I => \N__8067\
        );

    \I__838\ : InMux
    port map (
            O => \N__8070\,
            I => \N__8064\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__8067\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_3\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__8064\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_3\
        );

    \I__835\ : InMux
    port map (
            O => \N__8059\,
            I => \N__8056\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__8056\,
            I => \tx_fifo.lscc_fifo_inst.n5690\
        );

    \I__833\ : InMux
    port map (
            O => \N__8053\,
            I => \N__8050\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__8050\,
            I => \N__8046\
        );

    \I__831\ : InMux
    port map (
            O => \N__8049\,
            I => \N__8043\
        );

    \I__830\ : Span4Mux_h
    port map (
            O => \N__8046\,
            I => \N__8040\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__8043\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_6\
        );

    \I__828\ : Odrv4
    port map (
            O => \N__8040\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_6\
        );

    \I__827\ : CascadeMux
    port map (
            O => \N__8035\,
            I => \N__8031\
        );

    \I__826\ : InMux
    port map (
            O => \N__8034\,
            I => \N__8028\
        );

    \I__825\ : InMux
    port map (
            O => \N__8031\,
            I => \N__8025\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__8028\,
            I => \N__8022\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__8025\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_6\
        );

    \I__822\ : Odrv4
    port map (
            O => \N__8022\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_6\
        );

    \I__821\ : CascadeMux
    port map (
            O => \N__8017\,
            I => \tx_fifo.lscc_fifo_inst.n5696_cascade_\
        );

    \I__820\ : CascadeMux
    port map (
            O => \N__8014\,
            I => \N__8010\
        );

    \I__819\ : InMux
    port map (
            O => \N__8013\,
            I => \N__8007\
        );

    \I__818\ : InMux
    port map (
            O => \N__8010\,
            I => \N__8004\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__8007\,
            I => \N__8001\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__8004\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_6\
        );

    \I__815\ : Odrv4
    port map (
            O => \N__8001\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_6\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__7996\,
            I => \N__7993\
        );

    \I__813\ : InMux
    port map (
            O => \N__7993\,
            I => \N__7990\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__7990\,
            I => \N__7987\
        );

    \I__811\ : Odrv12
    port map (
            O => \N__7987\,
            I => \mem_LUT_data_raw_r_6\
        );

    \I__810\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7981\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__7981\,
            I => \tx_fifo.lscc_fifo_inst.n5702\
        );

    \I__808\ : CascadeMux
    port map (
            O => \N__7978\,
            I => \N__7975\
        );

    \I__807\ : InMux
    port map (
            O => \N__7975\,
            I => \N__7971\
        );

    \I__806\ : InMux
    port map (
            O => \N__7974\,
            I => \N__7968\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__7971\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_5\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__7968\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_5\
        );

    \I__803\ : CascadeMux
    port map (
            O => \N__7963\,
            I => \N__7960\
        );

    \I__802\ : InMux
    port map (
            O => \N__7960\,
            I => \N__7956\
        );

    \I__801\ : InMux
    port map (
            O => \N__7959\,
            I => \N__7953\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__7956\,
            I => \N__7950\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__7953\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_5\
        );

    \I__798\ : Odrv4
    port map (
            O => \N__7950\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_5\
        );

    \I__797\ : CascadeMux
    port map (
            O => \N__7945\,
            I => \N__7941\
        );

    \I__796\ : InMux
    port map (
            O => \N__7944\,
            I => \N__7938\
        );

    \I__795\ : InMux
    port map (
            O => \N__7941\,
            I => \N__7935\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__7938\,
            I => \N__7932\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__7935\,
            I => rx_shift_reg_6
        );

    \I__792\ : Odrv4
    port map (
            O => \N__7932\,
            I => rx_shift_reg_6
        );

    \I__791\ : CascadeMux
    port map (
            O => \N__7927\,
            I => \N__7924\
        );

    \I__790\ : InMux
    port map (
            O => \N__7924\,
            I => \N__7920\
        );

    \I__789\ : InMux
    port map (
            O => \N__7923\,
            I => \N__7917\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__7920\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_0\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__7917\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_0\
        );

    \I__786\ : InMux
    port map (
            O => \N__7912\,
            I => \N__7909\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__7909\,
            I => \tx_fifo.lscc_fifo_inst.n5666\
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__7906\,
            I => \N__7902\
        );

    \I__783\ : InMux
    port map (
            O => \N__7905\,
            I => \N__7899\
        );

    \I__782\ : InMux
    port map (
            O => \N__7902\,
            I => \N__7896\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__7899\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_0\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__7896\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_0\
        );

    \I__779\ : InMux
    port map (
            O => \N__7891\,
            I => \N__7885\
        );

    \I__778\ : InMux
    port map (
            O => \N__7890\,
            I => \N__7885\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__7885\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_2\
        );

    \I__776\ : CascadeMux
    port map (
            O => \N__7882\,
            I => \N__7878\
        );

    \I__775\ : InMux
    port map (
            O => \N__7881\,
            I => \N__7875\
        );

    \I__774\ : InMux
    port map (
            O => \N__7878\,
            I => \N__7872\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__7875\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_3\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__7872\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_3\
        );

    \I__771\ : InMux
    port map (
            O => \N__7867\,
            I => \N__7864\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__7864\,
            I => \N__7861\
        );

    \I__769\ : Span12Mux_h
    port map (
            O => \N__7861\,
            I => \N__7858\
        );

    \I__768\ : Span12Mux_v
    port map (
            O => \N__7858\,
            I => \N__7855\
        );

    \I__767\ : Odrv12
    port map (
            O => \N__7855\,
            I => \SOUT_c\
        );

    \I__766\ : InMux
    port map (
            O => \N__7852\,
            I => \N__7849\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__7849\,
            I => rx_shift_reg_0
        );

    \I__764\ : InMux
    port map (
            O => \N__7846\,
            I => \N__7843\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__7843\,
            I => \N__7840\
        );

    \I__762\ : Span12Mux_v
    port map (
            O => \N__7840\,
            I => \N__7837\
        );

    \I__761\ : Odrv12
    port map (
            O => \N__7837\,
            I => \FIFO_D28_c_28\
        );

    \I__760\ : IoInMux
    port map (
            O => \N__7834\,
            I => \N__7831\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__7831\,
            I => \N__7828\
        );

    \I__758\ : Span4Mux_s3_v
    port map (
            O => \N__7828\,
            I => \N__7825\
        );

    \I__757\ : Span4Mux_v
    port map (
            O => \N__7825\,
            I => \N__7822\
        );

    \I__756\ : Span4Mux_v
    port map (
            O => \N__7822\,
            I => \N__7819\
        );

    \I__755\ : Odrv4
    port map (
            O => \N__7819\,
            I => \DATA28_c_28\
        );

    \I__754\ : IoInMux
    port map (
            O => \N__7816\,
            I => \N__7813\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__7813\,
            I => \N__7810\
        );

    \I__752\ : Span4Mux_s1_v
    port map (
            O => \N__7810\,
            I => \N__7807\
        );

    \I__751\ : Sp12to4
    port map (
            O => \N__7807\,
            I => \N__7804\
        );

    \I__750\ : Span12Mux_s7_h
    port map (
            O => \N__7804\,
            I => \N__7801\
        );

    \I__749\ : Span12Mux_v
    port map (
            O => \N__7801\,
            I => \N__7798\
        );

    \I__748\ : Odrv12
    port map (
            O => \N__7798\,
            I => \SCK_c\
        );

    \I__747\ : InMux
    port map (
            O => \N__7795\,
            I => \N__7792\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__7792\,
            I => \N__7789\
        );

    \I__745\ : Span12Mux_v
    port map (
            O => \N__7789\,
            I => \N__7786\
        );

    \I__744\ : Odrv12
    port map (
            O => \N__7786\,
            I => \FIFO_D23_c_23\
        );

    \I__743\ : IoInMux
    port map (
            O => \N__7783\,
            I => \N__7780\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__7780\,
            I => \N__7777\
        );

    \I__741\ : Span4Mux_s3_v
    port map (
            O => \N__7777\,
            I => \N__7774\
        );

    \I__740\ : Span4Mux_h
    port map (
            O => \N__7774\,
            I => \N__7771\
        );

    \I__739\ : Sp12to4
    port map (
            O => \N__7771\,
            I => \N__7768\
        );

    \I__738\ : Span12Mux_h
    port map (
            O => \N__7768\,
            I => \N__7765\
        );

    \I__737\ : Odrv12
    port map (
            O => \N__7765\,
            I => \DATA23_c_23\
        );

    \I__736\ : CascadeMux
    port map (
            O => \N__7762\,
            I => \N__7757\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__7761\,
            I => \N__7753\
        );

    \I__734\ : InMux
    port map (
            O => \N__7760\,
            I => \N__7749\
        );

    \I__733\ : InMux
    port map (
            O => \N__7757\,
            I => \N__7746\
        );

    \I__732\ : InMux
    port map (
            O => \N__7756\,
            I => \N__7741\
        );

    \I__731\ : InMux
    port map (
            O => \N__7753\,
            I => \N__7741\
        );

    \I__730\ : InMux
    port map (
            O => \N__7752\,
            I => \N__7738\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__7749\,
            I => rx_buf_byte_0
        );

    \I__728\ : LocalMux
    port map (
            O => \N__7746\,
            I => rx_buf_byte_0
        );

    \I__727\ : LocalMux
    port map (
            O => \N__7741\,
            I => rx_buf_byte_0
        );

    \I__726\ : LocalMux
    port map (
            O => \N__7738\,
            I => rx_buf_byte_0
        );

    \I__725\ : InMux
    port map (
            O => \N__7729\,
            I => \N__7725\
        );

    \I__724\ : InMux
    port map (
            O => \N__7728\,
            I => \N__7722\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__7725\,
            I => \N__7719\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__7722\,
            I => rx_shift_reg_7
        );

    \I__721\ : Odrv4
    port map (
            O => \N__7719\,
            I => rx_shift_reg_7
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__7714\,
            I => \N__7711\
        );

    \I__719\ : InMux
    port map (
            O => \N__7711\,
            I => \N__7705\
        );

    \I__718\ : InMux
    port map (
            O => \N__7710\,
            I => \N__7705\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__7705\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_3\
        );

    \I__716\ : InMux
    port map (
            O => \N__7702\,
            I => \N__7699\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__7699\,
            I => \N__7696\
        );

    \I__714\ : Span4Mux_v
    port map (
            O => \N__7696\,
            I => \N__7693\
        );

    \I__713\ : Sp12to4
    port map (
            O => \N__7693\,
            I => \N__7690\
        );

    \I__712\ : Odrv12
    port map (
            O => \N__7690\,
            I => \FIFO_D31_c_31\
        );

    \I__711\ : IoInMux
    port map (
            O => \N__7687\,
            I => \N__7684\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__7684\,
            I => \N__7681\
        );

    \I__709\ : IoSpan4Mux
    port map (
            O => \N__7681\,
            I => \N__7678\
        );

    \I__708\ : Span4Mux_s2_v
    port map (
            O => \N__7678\,
            I => \N__7675\
        );

    \I__707\ : Sp12to4
    port map (
            O => \N__7675\,
            I => \N__7672\
        );

    \I__706\ : Span12Mux_v
    port map (
            O => \N__7672\,
            I => \N__7669\
        );

    \I__705\ : Odrv12
    port map (
            O => \N__7669\,
            I => \DATA31_c_31\
        );

    \I__704\ : InMux
    port map (
            O => \N__7666\,
            I => \N__7663\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__7663\,
            I => \N__7660\
        );

    \I__702\ : Span4Mux_h
    port map (
            O => \N__7660\,
            I => \N__7657\
        );

    \I__701\ : Span4Mux_v
    port map (
            O => \N__7657\,
            I => \N__7654\
        );

    \I__700\ : Span4Mux_v
    port map (
            O => \N__7654\,
            I => \N__7651\
        );

    \I__699\ : Odrv4
    port map (
            O => \N__7651\,
            I => \FIFO_D11_c_11\
        );

    \I__698\ : IoInMux
    port map (
            O => \N__7648\,
            I => \N__7645\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__7645\,
            I => \N__7642\
        );

    \I__696\ : IoSpan4Mux
    port map (
            O => \N__7642\,
            I => \N__7639\
        );

    \I__695\ : Span4Mux_s2_h
    port map (
            O => \N__7639\,
            I => \N__7636\
        );

    \I__694\ : Sp12to4
    port map (
            O => \N__7636\,
            I => \N__7633\
        );

    \I__693\ : Span12Mux_v
    port map (
            O => \N__7633\,
            I => \N__7630\
        );

    \I__692\ : Span12Mux_h
    port map (
            O => \N__7630\,
            I => \N__7627\
        );

    \I__691\ : Odrv12
    port map (
            O => \N__7627\,
            I => \DATA11_c_11\
        );

    \I__690\ : InMux
    port map (
            O => \N__7624\,
            I => \N__7620\
        );

    \I__689\ : InMux
    port map (
            O => \N__7623\,
            I => \N__7617\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__7620\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_0\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__7617\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_0\
        );

    \I__686\ : CascadeMux
    port map (
            O => \N__7612\,
            I => \N__7608\
        );

    \I__685\ : CascadeMux
    port map (
            O => \N__7611\,
            I => \N__7605\
        );

    \I__684\ : InMux
    port map (
            O => \N__7608\,
            I => \N__7602\
        );

    \I__683\ : InMux
    port map (
            O => \N__7605\,
            I => \N__7599\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__7602\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_0\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__7599\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_0\
        );

    \I__680\ : InMux
    port map (
            O => \N__7594\,
            I => \N__7591\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__7591\,
            I => rx_shift_reg_8
        );

    \I__678\ : IoInMux
    port map (
            O => \N__7588\,
            I => \N__7585\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__7585\,
            I => \N__7581\
        );

    \I__676\ : IoInMux
    port map (
            O => \N__7584\,
            I => \N__7578\
        );

    \I__675\ : IoSpan4Mux
    port map (
            O => \N__7581\,
            I => \N__7573\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__7578\,
            I => \N__7573\
        );

    \I__673\ : Span4Mux_s3_h
    port map (
            O => \N__7573\,
            I => \N__7570\
        );

    \I__672\ : Span4Mux_v
    port map (
            O => \N__7570\,
            I => \N__7567\
        );

    \I__671\ : Odrv4
    port map (
            O => \N__7567\,
            I => \FT_RD_c\
        );

    \I__670\ : InMux
    port map (
            O => \N__7564\,
            I => \N__7561\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__7561\,
            I => \N__7558\
        );

    \I__668\ : Sp12to4
    port map (
            O => \N__7558\,
            I => \N__7555\
        );

    \I__667\ : Span12Mux_v
    port map (
            O => \N__7555\,
            I => \N__7552\
        );

    \I__666\ : Odrv12
    port map (
            O => \N__7552\,
            I => \FIFO_D19_c_19\
        );

    \I__665\ : IoInMux
    port map (
            O => \N__7549\,
            I => \N__7546\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__7546\,
            I => \N__7543\
        );

    \I__663\ : Span4Mux_s3_v
    port map (
            O => \N__7543\,
            I => \N__7540\
        );

    \I__662\ : Span4Mux_v
    port map (
            O => \N__7540\,
            I => \N__7537\
        );

    \I__661\ : Sp12to4
    port map (
            O => \N__7537\,
            I => \N__7534\
        );

    \I__660\ : Span12Mux_h
    port map (
            O => \N__7534\,
            I => \N__7531\
        );

    \I__659\ : Span12Mux_v
    port map (
            O => \N__7531\,
            I => \N__7528\
        );

    \I__658\ : Odrv12
    port map (
            O => \N__7528\,
            I => \DATA19_c_19\
        );

    \I__657\ : InMux
    port map (
            O => \N__7525\,
            I => \N__7522\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__7522\,
            I => \N__7519\
        );

    \I__655\ : Span4Mux_v
    port map (
            O => \N__7519\,
            I => \N__7516\
        );

    \I__654\ : Sp12to4
    port map (
            O => \N__7516\,
            I => \N__7513\
        );

    \I__653\ : Span12Mux_h
    port map (
            O => \N__7513\,
            I => \N__7510\
        );

    \I__652\ : Span12Mux_v
    port map (
            O => \N__7510\,
            I => \N__7507\
        );

    \I__651\ : Odrv12
    port map (
            O => \N__7507\,
            I => \FIFO_D14_c_14\
        );

    \I__650\ : IoInMux
    port map (
            O => \N__7504\,
            I => \N__7501\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__7501\,
            I => \N__7498\
        );

    \I__648\ : IoSpan4Mux
    port map (
            O => \N__7498\,
            I => \N__7495\
        );

    \I__647\ : Span4Mux_s3_h
    port map (
            O => \N__7495\,
            I => \N__7492\
        );

    \I__646\ : Sp12to4
    port map (
            O => \N__7492\,
            I => \N__7489\
        );

    \I__645\ : Span12Mux_s11_h
    port map (
            O => \N__7489\,
            I => \N__7486\
        );

    \I__644\ : Span12Mux_h
    port map (
            O => \N__7486\,
            I => \N__7483\
        );

    \I__643\ : Odrv12
    port map (
            O => \N__7483\,
            I => \DATA14_c_14\
        );

    \I__642\ : InMux
    port map (
            O => \N__7480\,
            I => \N__7477\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__7477\,
            I => \N__7474\
        );

    \I__640\ : Span4Mux_v
    port map (
            O => \N__7474\,
            I => \N__7471\
        );

    \I__639\ : Sp12to4
    port map (
            O => \N__7471\,
            I => \N__7468\
        );

    \I__638\ : Odrv12
    port map (
            O => \N__7468\,
            I => \FIFO_D30_c_30\
        );

    \I__637\ : IoInMux
    port map (
            O => \N__7465\,
            I => \N__7462\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__7462\,
            I => \N__7459\
        );

    \I__635\ : Span4Mux_s1_v
    port map (
            O => \N__7459\,
            I => \N__7456\
        );

    \I__634\ : Span4Mux_v
    port map (
            O => \N__7456\,
            I => \N__7453\
        );

    \I__633\ : Span4Mux_v
    port map (
            O => \N__7453\,
            I => \N__7450\
        );

    \I__632\ : Span4Mux_v
    port map (
            O => \N__7450\,
            I => \N__7447\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__7447\,
            I => \DATA30_c_30\
        );

    \INVspi0.tx_shift_reg_i0C\ : INV
    port map (
            O => \INVspi0.tx_shift_reg_i0C_net\,
            I => \N__10125\
        );

    \INVspi0.tx_shift_reg_i15C\ : INV
    port map (
            O => \INVspi0.tx_shift_reg_i15C_net\,
            I => \N__10123\
        );

    \INVspi0.tx_shift_reg_i6C\ : INV
    port map (
            O => \INVspi0.tx_shift_reg_i6C_net\,
            I => \N__10119\
        );

    \INVspi0.tx_shift_reg_i8C\ : INV
    port map (
            O => \INVspi0.tx_shift_reg_i8C_net\,
            I => \N__10107\
        );

    \IN_MUX_bfv_16_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_5_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pc_tx.n4872\,
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_13_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_6_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pc_rx.n4814\,
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_23_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_23_5_0_\
        );

    \IN_MUX_bfv_23_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n4830,
            carryinitout => \bfn_23_6_0_\
        );

    \IN_MUX_bfv_23_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n4838,
            carryinitout => \bfn_23_7_0_\
        );

    \IN_MUX_bfv_23_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n4846,
            carryinitout => \bfn_23_8_0_\
        );

    \IN_MUX_bfv_17_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_8_0_\
        );

    \IN_MUX_bfv_17_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_7_0_\
        );

    \IN_MUX_bfv_15_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_8_0_\
        );

    \IN_MUX_bfv_15_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \bluejay_data_inst.n4854\,
            carryinitout => \bfn_15_9_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i1_2_lut_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__18667\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19507\,
            lcout => \FT_RD_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2715_2_lut_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7564\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18958\,
            lcout => \DATA19_c_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2722_2_lut_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7525\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18955\,
            lcout => \DATA14_c_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2702_2_lut_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18957\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7480\,
            lcout => \DATA30_c_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2701_2_lut_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7702\,
            in2 => \_gnd_net_\,
            in3 => \N__18956\,
            lcout => \DATA31_c_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i38_39_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__12169\,
            in1 => \N__10699\,
            in2 => \N__7762\,
            in3 => \N__7905\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i230_231_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__7624\,
            in1 => \N__10698\,
            in2 => \N__7761\,
            in3 => \N__12170\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i326_327_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__12168\,
            in1 => \N__7756\,
            in2 => \N__7612\,
            in3 => \N__10572\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2725_2_lut_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18970\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7666\,
            lcout => \DATA11_c_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i7_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8701\,
            in1 => \N__7594\,
            in2 => \_gnd_net_\,
            in3 => \N__10262\,
            lcout => rx_buf_byte_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i0_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8257\,
            in1 => \N__7752\,
            in2 => \_gnd_net_\,
            in3 => \N__8700\,
            lcout => rx_buf_byte_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_4713_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__7623\,
            in1 => \N__12400\,
            in2 => \N__7611\,
            in3 => \N__14261\,
            lcout => \tx_fifo.lscc_fifo_inst.n5666\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__3_i9_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7729\,
            in2 => \_gnd_net_\,
            in3 => \N__11185\,
            lcout => rx_shift_reg_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i248_249_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__8049\,
            in1 => \N__10728\,
            in2 => \N__8586\,
            in3 => \N__12186\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__3_i8_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7944\,
            in2 => \_gnd_net_\,
            in3 => \N__11181\,
            lcout => rx_shift_reg_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i6_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7728\,
            in1 => \N__8577\,
            in2 => \_gnd_net_\,
            in3 => \N__8699\,
            lcout => rx_buf_byte_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i341_342_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__8100\,
            in1 => \N__12106\,
            in2 => \N__10624\,
            in3 => \N__8335\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i239_240_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__10733\,
            in1 => \N__8285\,
            in2 => \N__7714\,
            in3 => \N__12107\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_4733_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__14258\,
            in1 => \N__7710\,
            in2 => \N__7882\,
            in3 => \N__12403\,
            lcout => \tx_fifo.lscc_fifo_inst.n5690\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i245_246_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__10734\,
            in1 => \N__8334\,
            in2 => \N__8119\,
            in3 => \N__12108\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i47_48_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__12105\,
            in1 => \N__8086\,
            in2 => \N__8290\,
            in3 => \N__10735\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i53_54_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__12181\,
            in1 => \N__7959\,
            in2 => \N__10741\,
            in3 => \N__8328\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i149_150_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__10617\,
            in1 => \N__8327\,
            in2 => \N__7978\,
            in3 => \N__12182\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__3_i2_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11177\,
            in2 => \_gnd_net_\,
            in3 => \N__7852\,
            lcout => rx_shift_reg_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10075\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__3_i1_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__7867\,
            in1 => \N__11176\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => rx_shift_reg_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10075\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__3_i7_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__11180\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8712\,
            lcout => rx_shift_reg_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10075\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__3_i5_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11178\,
            in2 => \_gnd_net_\,
            in3 => \N__8232\,
            lcout => rx_shift_reg_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10075\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__3_i6_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__11179\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8301\,
            lcout => rx_shift_reg_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10075\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2704_2_lut_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7846\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18960\,
            lcout => \DATA28_c_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i2_3_lut_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__14475\,
            in1 => \N__10026\,
            in2 => \_gnd_net_\,
            in3 => \N__8205\,
            lcout => \SCK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2709_2_lut_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7795\,
            in2 => \_gnd_net_\,
            in3 => \N__18969\,
            lcout => \DATA23_c_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i134_135_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__7760\,
            in1 => \N__10571\,
            in2 => \N__7927\,
            in3 => \N__12171\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i1_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__7923\,
            in1 => \N__7912\,
            in2 => \N__7906\,
            in3 => \N__12401\,
            lcout => \mem_LUT_data_raw_r_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19337\,
            ce => \N__11338\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i44_45_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__8347\,
            in1 => \N__10723\,
            in2 => \N__12188\,
            in3 => \N__8445\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_4708_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__7890\,
            in1 => \N__12382\,
            in2 => \N__8412\,
            in3 => \N__14259\,
            lcout => \tx_fifo.lscc_fifo_inst.n5660\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i236_237_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__7891\,
            in1 => \N__10722\,
            in2 => \N__12187\,
            in3 => \N__8444\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i6_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__8388\,
            in1 => \N__11899\,
            in2 => \N__7996\,
            in3 => \N__16576\,
            lcout => fifo_temp_output_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.t_FSM_i5_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__9490\,
            in1 => \N__12969\,
            in2 => \N__9589\,
            in3 => \N__9433\,
            lcout => \spi0.n490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10118\,
            ce => 'H',
            sr => \N__16544\
        );

    \tx_fifo.lscc_fifo_inst.i152_153_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__10613\,
            in1 => \N__8581\,
            in2 => \N__8014\,
            in3 => \N__12160\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i140_141_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__12158\,
            in1 => \N__8443\,
            in2 => \N__8373\,
            in3 => \N__10615\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i143_144_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__10612\,
            in1 => \N__8073\,
            in2 => \N__12190\,
            in3 => \N__8281\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i335_336_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__12159\,
            in1 => \N__7881\,
            in2 => \N__8289\,
            in3 => \N__10616\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i329_330_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__10614\,
            in1 => \N__8514\,
            in2 => \N__9322\,
            in3 => \N__12161\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i56_57_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__8582\,
            in1 => \N__10729\,
            in2 => \N__8035\,
            in3 => \N__12162\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__8118\,
            in1 => \N__12399\,
            in2 => \N__8101\,
            in3 => \N__14257\,
            lcout => \tx_fifo.lscc_fifo_inst.n5702\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i8_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100110101000"
        )
    port map (
            in0 => \N__9691\,
            in1 => \N__12381\,
            in2 => \N__8755\,
            in3 => \N__8769\,
            lcout => \mem_LUT_data_raw_r_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19326\,
            ce => \N__11330\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i4_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__12378\,
            in1 => \N__8085\,
            in2 => \N__8074\,
            in3 => \N__8059\,
            lcout => \mem_LUT_data_raw_r_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19326\,
            ce => \N__11330\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_4738_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__8053\,
            in1 => \N__12377\,
            in2 => \N__8551\,
            in3 => \N__14260\,
            lcout => OPEN,
            ltout => \tx_fifo.lscc_fifo_inst.n5696_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i7_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__12379\,
            in1 => \N__8034\,
            in2 => \N__8017\,
            in3 => \N__8013\,
            lcout => \mem_LUT_data_raw_r_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19326\,
            ce => \N__11330\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i6_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__7984\,
            in1 => \N__7974\,
            in2 => \N__7963\,
            in3 => \N__12380\,
            lcout => \mem_LUT_data_raw_r_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19326\,
            ce => \N__11330\,
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i5_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__8684\,
            in1 => \_gnd_net_\,
            in2 => \N__7945\,
            in3 => \N__8326\,
            lcout => rx_buf_byte_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i1_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8242\,
            in1 => \N__9301\,
            in2 => \_gnd_net_\,
            in3 => \N__8681\,
            lcout => rx_buf_byte_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__3_i4_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8241\,
            in2 => \_gnd_net_\,
            in3 => \N__11169\,
            lcout => rx_shift_reg_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i3_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8305\,
            in1 => \N__8270\,
            in2 => \_gnd_net_\,
            in3 => \N__8683\,
            lcout => rx_buf_byte_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__3_i3_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8253\,
            in2 => \_gnd_net_\,
            in3 => \N__11168\,
            lcout => rx_shift_reg_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i2_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8233\,
            in1 => \N__8431\,
            in2 => \_gnd_net_\,
            in3 => \N__8682\,
            lcout => rx_buf_byte_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.CS_81_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9916\,
            lcout => \SEN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10082\,
            ce => 'H',
            sr => \N__16545\
        );

    \bluejay_data_inst.i2707_2_lut_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18962\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8194\,
            lcout => \DATA25_c_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2703_2_lut_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8152\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18961\,
            lcout => \DATA29_c_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Bit_Index_i2_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9166\,
            in1 => \N__9136\,
            in2 => \_gnd_net_\,
            in3 => \N__9066\,
            lcout => \pc_tx.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19347\,
            ce => \N__9850\,
            sr => \N__9085\
        );

    \pc_tx.r_Bit_Index_i1_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__9067\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9165\,
            lcout => \pc_tx.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19347\,
            ce => \N__9850\,
            sr => \N__9085\
        );

    \tx_fifo.lscc_fifo_inst.i332_333_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__12167\,
            in1 => \N__8449\,
            in2 => \N__8413\,
            in3 => \N__10599\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i41_42_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__10701\,
            in1 => \N__8500\,
            in2 => \N__12189\,
            in3 => \N__9327\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i233_234_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__12166\,
            in1 => \N__8535\,
            in2 => \N__9328\,
            in3 => \N__10700\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i6_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9241\,
            in1 => \N__8395\,
            in2 => \_gnd_net_\,
            in3 => \N__9178\,
            lcout => \r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i4_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__16575\,
            in1 => \N__8997\,
            in2 => \N__8482\,
            in3 => \N__11901\,
            lcout => fifo_temp_output_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2_2_lut_3_lut_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9134\,
            in1 => \N__9164\,
            in2 => \_gnd_net_\,
            in3 => \N__9064\,
            lcout => \pc_tx.n3763\,
            ltout => \pc_tx.n3763_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Bit_Index_i0_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010010101010"
        )
    port map (
            in0 => \N__9065\,
            in1 => \N__15536\,
            in2 => \N__8377\,
            in3 => \N__9846\,
            lcout => \pc_tx.r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i3_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101111001000"
        )
    port map (
            in0 => \N__8374\,
            in1 => \N__8353\,
            in2 => \N__12402\,
            in3 => \N__8346\,
            lcout => \mem_LUT_data_raw_r_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19338\,
            ce => \N__11334\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_4718_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__8536\,
            in1 => \N__12389\,
            in2 => \N__8521\,
            in3 => \N__14266\,
            lcout => OPEN,
            ltout => \tx_fifo.lscc_fifo_inst.n5672_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i2_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__12391\,
            in1 => \N__8499\,
            in2 => \N__8488\,
            in3 => \N__9279\,
            lcout => \mem_LUT_data_raw_r_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19338\,
            ce => \N__11334\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_4723_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000111000"
        )
    port map (
            in0 => \N__10150\,
            in1 => \N__12390\,
            in2 => \N__14265\,
            in3 => \N__9021\,
            lcout => OPEN,
            ltout => \tx_fifo.lscc_fifo_inst.n5678_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i5_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__12392\,
            in1 => \N__9198\,
            in2 => \N__8485\,
            in3 => \N__8736\,
            lcout => \mem_LUT_data_raw_r_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19338\,
            ce => \N__11334\,
            sr => \_gnd_net_\
        );

    \spi0.t_FSM_i15_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000100"
        )
    port map (
            in0 => \N__12944\,
            in1 => \N__8464\,
            in2 => \N__9520\,
            in3 => \N__9423\,
            lcout => \spi0.n480\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10126\,
            ce => 'H',
            sr => \N__16565\
        );

    \spi0.mux_473_i2_4_lut_4_lut_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__13043\,
            in1 => \N__9784\,
            in2 => \N__9540\,
            in3 => \N__12937\,
            lcout => \spi0.state_next_1\,
            ltout => \spi0.state_next_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.t_FSM_i0_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111011110"
        )
    port map (
            in0 => \N__12938\,
            in1 => \N__8473\,
            in2 => \N__8467\,
            in3 => \N__9417\,
            lcout => \spi0.n495\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10126\,
            ce => 'H',
            sr => \N__16565\
        );

    \spi0.t_FSM_i14_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000010000"
        )
    port map (
            in0 => \N__9422\,
            in1 => \N__9504\,
            in2 => \N__8458\,
            in3 => \N__12943\,
            lcout => \spi0.n481\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10126\,
            ce => 'H',
            sr => \N__16565\
        );

    \spi0.t_FSM_i13_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000100"
        )
    port map (
            in0 => \N__12942\,
            in1 => \N__8647\,
            in2 => \N__9519\,
            in3 => \N__9421\,
            lcout => \spi0.n482\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10126\,
            ce => 'H',
            sr => \N__16565\
        );

    \spi0.t_FSM_i12_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000010000"
        )
    port map (
            in0 => \N__9420\,
            in1 => \N__9503\,
            in2 => \N__8641\,
            in3 => \N__12941\,
            lcout => \spi0.n483\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10126\,
            ce => 'H',
            sr => \N__16565\
        );

    \spi0.t_FSM_i11_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000100"
        )
    port map (
            in0 => \N__12940\,
            in1 => \N__8632\,
            in2 => \N__9518\,
            in3 => \N__9419\,
            lcout => \spi0.n484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10126\,
            ce => 'H',
            sr => \N__16565\
        );

    \spi0.t_FSM_i10_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000010000"
        )
    port map (
            in0 => \N__9418\,
            in1 => \N__9502\,
            in2 => \N__8602\,
            in3 => \N__12939\,
            lcout => \spi0.n485\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10126\,
            ce => 'H',
            sr => \N__16565\
        );

    \spi0.t_FSM_i6_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__12930\,
            in1 => \N__9491\,
            in2 => \N__8626\,
            in3 => \N__9429\,
            lcout => \state_next_2__N_454\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10111\,
            ce => 'H',
            sr => \N__16578\
        );

    \spi0.i1_2_lut_3_lut_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__9571\,
            in1 => \N__11726\,
            in2 => \_gnd_net_\,
            in3 => \N__12929\,
            lcout => \spi0.n1005\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.t_FSM_i7_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__12931\,
            in1 => \N__9492\,
            in2 => \N__9577\,
            in3 => \N__9430\,
            lcout => \spi0.n488\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10111\,
            ce => 'H',
            sr => \N__16578\
        );

    \spi0.t_FSM_i8_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000100"
        )
    port map (
            in0 => \N__9431\,
            in1 => \N__8617\,
            in2 => \N__9515\,
            in3 => \N__12932\,
            lcout => \spi0.n487\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10111\,
            ce => 'H',
            sr => \N__16578\
        );

    \spi0.t_FSM_i9_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__12933\,
            in1 => \N__9493\,
            in2 => \N__8611\,
            in3 => \N__9432\,
            lcout => \spi0.n486\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10111\,
            ce => 'H',
            sr => \N__16578\
        );

    \tx_fifo.lscc_fifo_inst.i344_345_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__8550\,
            in1 => \N__10605\,
            in2 => \N__8593\,
            in3 => \N__12153\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i347_348_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__12151\,
            in1 => \N__10283\,
            in2 => \N__10623\,
            in3 => \N__9705\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i59_60_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__10740\,
            in1 => \N__10284\,
            in2 => \N__8770\,
            in3 => \N__12154\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i155_156_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__12150\,
            in1 => \N__8754\,
            in2 => \N__10622\,
            in3 => \N__10282\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.state_reg_2__I_0_108_i5_3_lut_3_lut_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__13053\,
            in1 => \N__12945\,
            in2 => \_gnd_net_\,
            in3 => \N__11736\,
            lcout => \rx_shift_reg_15__N_461\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i146_147_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__10172\,
            in1 => \N__10604\,
            in2 => \N__8737\,
            in3 => \N__12152\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i6_4_lut_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__8850\,
            in1 => \N__8916\,
            in2 => \N__8815\,
            in3 => \N__8883\,
            lcout => OPEN,
            ltout => \spi0.n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i4676_4_lut_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8832\,
            in1 => \N__8932\,
            in2 => \N__8719\,
            in3 => \N__8653\,
            lcout => \spi0.n2715\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i4_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8716\,
            in1 => \N__10171\,
            in2 => \_gnd_net_\,
            in3 => \N__8680\,
            lcout => rx_buf_byte_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10096\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i2_2_lut_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8865\,
            in2 => \_gnd_net_\,
            in3 => \N__8898\,
            lcout => \spi0.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.spi_clk_counter_701__i0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8931\,
            in2 => \_gnd_net_\,
            in3 => \N__8920\,
            lcout => \spi0.spi_clk_counter_0\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \spi0.n4874\,
            clk => \N__19334\,
            ce => 'H',
            sr => \N__9901\
        );

    \spi0.spi_clk_counter_701__i1_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8917\,
            in2 => \N__17112\,
            in3 => \N__8905\,
            lcout => \spi0.spi_clk_counter_1\,
            ltout => OPEN,
            carryin => \spi0.n4874\,
            carryout => \spi0.n4875\,
            clk => \N__19334\,
            ce => 'H',
            sr => \N__9901\
        );

    \spi0.spi_clk_counter_701__i2_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17096\,
            in2 => \N__8902\,
            in3 => \N__8887\,
            lcout => \spi0.spi_clk_counter_2\,
            ltout => OPEN,
            carryin => \spi0.n4875\,
            carryout => \spi0.n4876\,
            clk => \N__19334\,
            ce => 'H',
            sr => \N__9901\
        );

    \spi0.spi_clk_counter_701__i3_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8884\,
            in2 => \N__17113\,
            in3 => \N__8872\,
            lcout => \spi0.spi_clk_counter_3\,
            ltout => OPEN,
            carryin => \spi0.n4876\,
            carryout => \spi0.n4877\,
            clk => \N__19334\,
            ce => 'H',
            sr => \N__9901\
        );

    \spi0.spi_clk_counter_701__i4_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17100\,
            in2 => \N__8869\,
            in3 => \N__8854\,
            lcout => \spi0.spi_clk_counter_4\,
            ltout => OPEN,
            carryin => \spi0.n4877\,
            carryout => \spi0.n4878\,
            clk => \N__19334\,
            ce => 'H',
            sr => \N__9901\
        );

    \spi0.spi_clk_counter_701__i5_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8851\,
            in2 => \N__17114\,
            in3 => \N__8839\,
            lcout => \spi0.spi_clk_counter_5\,
            ltout => OPEN,
            carryin => \spi0.n4878\,
            carryout => \spi0.n4879\,
            clk => \N__19334\,
            ce => 'H',
            sr => \N__9901\
        );

    \spi0.spi_clk_counter_701__i6_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17104\,
            in2 => \N__8836\,
            in3 => \N__8821\,
            lcout => \spi0.spi_clk_counter_6\,
            ltout => OPEN,
            carryin => \spi0.n4879\,
            carryout => \spi0.n4880\,
            clk => \N__19334\,
            ce => 'H',
            sr => \N__9901\
        );

    \spi0.spi_clk_counter_701__i7_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17105\,
            in1 => \N__8814\,
            in2 => \_gnd_net_\,
            in3 => \N__8818\,
            lcout => \spi0.spi_clk_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19334\,
            ce => 'H',
            sr => \N__9901\
        );

    \bluejay_data_inst.i2716_2_lut_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8800\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18959\,
            lcout => \DATA18_c_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i5_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8956\,
            in1 => \N__9724\,
            in2 => \_gnd_net_\,
            in3 => \N__9240\,
            lcout => \r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19352\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i2_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__8986\,
            in1 => \N__11900\,
            in2 => \N__9010\,
            in3 => \N__16574\,
            lcout => fifo_temp_output_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19352\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Active_46_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111110000"
        )
    port map (
            in0 => \N__15523\,
            in1 => \N__16178\,
            in2 => \N__10994\,
            in3 => \N__8938\,
            lcout => tx_uart_active_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19352\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i3_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9358\,
            in1 => \N__9238\,
            in2 => \_gnd_net_\,
            in3 => \N__8974\,
            lcout => \r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19352\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i4_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8947\,
            in1 => \N__8998\,
            in2 => \_gnd_net_\,
            in3 => \N__9239\,
            lcout => \r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19352\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i2_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8965\,
            in1 => \N__8985\,
            in2 => \_gnd_net_\,
            in3 => \N__9237\,
            lcout => \r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19352\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i4551_3_lut_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8973\,
            in1 => \N__8964\,
            in2 => \_gnd_net_\,
            in3 => \N__9061\,
            lcout => \pc_tx.n5509\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i4553_3_lut_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9060\,
            in1 => \N__8955\,
            in2 => \_gnd_net_\,
            in3 => \N__8946\,
            lcout => \pc_tx.n5511\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i4645_4_lut_4_lut_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100000010000"
        )
    port map (
            in0 => \N__15526\,
            in1 => \N__15579\,
            in2 => \N__10237\,
            in3 => \N__15454\,
            lcout => n5414,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i4554_3_lut_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9075\,
            in1 => \N__9177\,
            in2 => \_gnd_net_\,
            in3 => \N__9062\,
            lcout => OPEN,
            ltout => \pc_tx.n5512_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Bit_Index_1__bdd_4_lut_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__9133\,
            in1 => \N__9163\,
            in2 => \N__9145\,
            in3 => \N__9142\,
            lcout => OPEN,
            ltout => \pc_tx.n5654_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.n5654_bdd_4_lut_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__9135\,
            in1 => \N__9028\,
            in2 => \N__9112\,
            in3 => \N__9109\,
            lcout => OPEN,
            ltout => \pc_tx.o_Tx_Serial_N_354_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_SM_Main_2__I_0_55_i3_3_lut_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15518\,
            in2 => \N__9103\,
            in3 => \N__15580\,
            lcout => \pc_tx.n3_adj_632\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i4680_2_lut_3_lut_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__15517\,
            in1 => \N__9871\,
            in2 => \_gnd_net_\,
            in3 => \N__9839\,
            lcout => \pc_tx.n5486\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2_3_lut_4_lut_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__15525\,
            in1 => \N__16152\,
            in2 => \N__10236\,
            in3 => \N__15578\,
            lcout => n2366,
            ltout => \n2366_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i7_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__9076\,
            in1 => \_gnd_net_\,
            in2 => \N__9079\,
            in3 => \N__11275\,
            lcout => \r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i4550_3_lut_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9264\,
            in1 => \N__9207\,
            in2 => \_gnd_net_\,
            in3 => \N__9063\,
            lcout => \pc_tx.n5508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i338_339_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__12163\,
            in1 => \N__10193\,
            in2 => \N__10621\,
            in3 => \N__9022\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i3_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__16547\,
            in1 => \N__9370\,
            in2 => \N__11902\,
            in3 => \N__9354\,
            lcout => fifo_temp_output_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i0_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__9255\,
            in1 => \N__11895\,
            in2 => \N__9343\,
            in3 => \N__16546\,
            lcout => fifo_temp_output_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i137_138_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__9323\,
            in1 => \N__10600\,
            in2 => \N__9280\,
            in3 => \N__12165\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i1_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__9236\,
            in1 => \_gnd_net_\,
            in2 => \N__9670\,
            in3 => \N__9265\,
            lcout => \r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i0_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9256\,
            in1 => \N__9235\,
            in2 => \_gnd_net_\,
            in3 => \N__9208\,
            lcout => \r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i50_51_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__12164\,
            in1 => \N__9199\,
            in2 => \N__10198\,
            in3 => \N__10721\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i1230_2_lut_4_lut_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100000000"
        )
    port map (
            in0 => \N__11721\,
            in1 => \N__12925\,
            in2 => \N__9575\,
            in3 => \N__13036\,
            lcout => \spi0.n2120\,
            ltout => \spi0.n2120_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.state_reg_i2_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001111100010"
        )
    port map (
            in0 => \N__13039\,
            in1 => \N__9783\,
            in2 => \N__9187\,
            in3 => \N__9184\,
            lcout => state_reg_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10113\,
            ce => 'H',
            sr => \N__16543\
        );

    \spi0.i4644_2_lut_3_lut_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__11722\,
            in1 => \N__12926\,
            in2 => \_gnd_net_\,
            in3 => \N__9816\,
            lcout => \spi0.n5552\,
            ltout => \spi0.n5552_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.mux_473_i3_4_lut_4_lut_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000110010"
        )
    port map (
            in0 => \N__13037\,
            in1 => \N__9781\,
            in2 => \N__9607\,
            in3 => \N__9755\,
            lcout => OPEN,
            ltout => \spi0.state_next_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i1_4_lut_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__11723\,
            in1 => \N__13038\,
            in2 => \N__9604\,
            in3 => \N__9739\,
            lcout => \spi0.n4\,
            ltout => \spi0.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.t_FSM_i3_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100100000000"
        )
    port map (
            in0 => \N__12927\,
            in1 => \N__9516\,
            in2 => \N__9601\,
            in3 => \N__9817\,
            lcout => \spi0.n492\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10113\,
            ce => 'H',
            sr => \N__16543\
        );

    \spi0.state_reg_i0_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__9782\,
            in1 => \_gnd_net_\,
            in2 => \N__9760\,
            in3 => \N__9790\,
            lcout => state_reg_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10113\,
            ce => 'H',
            sr => \N__16543\
        );

    \spi0.t_FSM_i4_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__12928\,
            in1 => \N__9517\,
            in2 => \N__9598\,
            in3 => \N__9416\,
            lcout => \spi0.n491\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10113\,
            ce => 'H',
            sr => \N__16543\
        );

    \i490_4_lut_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__13031\,
            in1 => \N__11725\,
            in2 => \N__9576\,
            in3 => \N__12919\,
            lcout => n982,
            ltout => \n982_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.state_reg_i1_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__12920\,
            in1 => \N__9541\,
            in2 => \N__9523\,
            in3 => \N__13033\,
            lcout => state_reg_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10083\,
            ce => 'H',
            sr => \N__16523\
        );

    \spi0.t_FSM_i2_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100000000"
        )
    port map (
            in0 => \N__9425\,
            in1 => \N__12922\,
            in2 => \N__9514\,
            in3 => \N__9826\,
            lcout => \spi0.state_next_2__N_452\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10083\,
            ce => 'H',
            sr => \N__16523\
        );

    \spi0.t_FSM_i1_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__12921\,
            in1 => \N__9486\,
            in2 => \N__9442\,
            in3 => \N__9424\,
            lcout => \spi0.state_next_2__N_453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10083\,
            ce => 'H',
            sr => \N__16523\
        );

    \spi0.i29_3_lut_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14446\,
            in1 => \N__12917\,
            in2 => \_gnd_net_\,
            in3 => \N__9825\,
            lcout => \spi0.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i4639_3_lut_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__12918\,
            in1 => \N__13030\,
            in2 => \_gnd_net_\,
            in3 => \N__9815\,
            lcout => OPEN,
            ltout => \spi0.n5561_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i28_4_lut_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011110011"
        )
    port map (
            in0 => \N__13032\,
            in1 => \N__11724\,
            in2 => \N__9799\,
            in3 => \N__9796\,
            lcout => \spi0.n13\,
            ltout => \spi0.n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.mux_473_i1_3_lut_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001101"
        )
    port map (
            in0 => \N__9780\,
            in1 => \N__9759\,
            in2 => \N__9742\,
            in3 => \_gnd_net_\,
            lcout => \spi0.state_next_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i5_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__16413\,
            in1 => \N__9733\,
            in2 => \N__11894\,
            in3 => \N__9717\,
            lcout => fifo_temp_output_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_4728_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__10248\,
            in1 => \N__12370\,
            in2 => \N__9706\,
            in3 => \N__14233\,
            lcout => \tx_fifo.lscc_fifo_inst.n5684\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__9663\,
            in1 => \N__11876\,
            in2 => \N__9682\,
            in3 => \N__16412\,
            lcout => fifo_temp_output_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2728_2_lut_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18881\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9652\,
            lcout => \DATA8_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.CS_w_79_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11737\,
            in2 => \_gnd_net_\,
            in3 => \N__13054\,
            lcout => \spi0.CS_w\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10025\,
            ce => 'H',
            sr => \N__12970\
        );

    \spi0.spi_clk_76_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__9978\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9897\,
            lcout => \spi0.spi_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_SM_Main_i1_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__15522\,
            in1 => \N__15585\,
            in2 => \_gnd_net_\,
            in3 => \N__15459\,
            lcout => \r_SM_Main_1_adj_660\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19357\,
            ce => 'H',
            sr => \N__16179\
        );

    \pc_tx.i1_3_lut_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__10485\,
            in1 => \N__10965\,
            in2 => \_gnd_net_\,
            in3 => \N__10500\,
            lcout => OPEN,
            ltout => \pc_tx.n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2_4_lut_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__10920\,
            in1 => \N__10935\,
            in2 => \N__9880\,
            in3 => \N__10132\,
            lcout => OPEN,
            ltout => \pc_tx.n4905_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2_4_lut_adj_26_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__10890\,
            in1 => \N__10905\,
            in2 => \N__9877\,
            in3 => \N__10872\,
            lcout => \pc_tx.r_SM_Main_2_N_322_1\,
            ltout => \pc_tx.r_SM_Main_2_N_322_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_SM_Main_i0_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15577\,
            in2 => \N__9874\,
            in3 => \N__9856\,
            lcout => \pc_tx.r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19353\,
            ce => 'H',
            sr => \N__16180\
        );

    \pc_tx.i1179_4_lut_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__15453\,
            in1 => \N__15505\,
            in2 => \N__10235\,
            in3 => \N__9870\,
            lcout => \pc_tx.n2069\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i1_3_lut_4_lut_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__16151\,
            in1 => \N__15576\,
            in2 => \N__15524\,
            in3 => \N__15452\,
            lcout => \pc_tx.n5484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2_2_lut_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10950\,
            in2 => \_gnd_net_\,
            in3 => \N__10470\,
            lcout => \pc_tx.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.state_reg_2__I_0_101_i5_2_lut_3_lut_3_lut_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__11734\,
            in1 => \N__13051\,
            in2 => \_gnd_net_\,
            in3 => \N__12961\,
            lcout => n5_adj_667,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i4684_4_lut_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000001"
        )
    port map (
            in0 => \N__15581\,
            in1 => \N__16177\,
            in2 => \N__15540\,
            in3 => \N__15455\,
            lcout => \pc_tx.n2739\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.busy_86_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__11733\,
            in1 => \N__13050\,
            in2 => \_gnd_net_\,
            in3 => \N__12960\,
            lcout => spi_busy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i8_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__11132\,
            in1 => \N__13705\,
            in2 => \N__11079\,
            in3 => \N__10294\,
            lcout => tx_shift_reg_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i8C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i4_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__9922\,
            in1 => \N__11130\,
            in2 => \N__12478\,
            in3 => \N__11057\,
            lcout => tx_shift_reg_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i8C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i1_2_lut_3_lut_adj_63_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__11717\,
            in1 => \N__13035\,
            in2 => \_gnd_net_\,
            in3 => \N__12924\,
            lcout => n2446,
            ltout => \n2446_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i5_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__12439\,
            in1 => \N__11131\,
            in2 => \N__9937\,
            in3 => \N__9934\,
            lcout => tx_shift_reg_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i8C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i9_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__11133\,
            in1 => \N__11419\,
            in2 => \N__11080\,
            in3 => \N__9928\,
            lcout => tx_shift_reg_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i8C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i3_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__11209\,
            in1 => \N__11129\,
            in2 => \N__13777\,
            in3 => \N__11056\,
            lcout => tx_shift_reg_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i8C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i11_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__11128\,
            in1 => \N__13747\,
            in2 => \N__11078\,
            in3 => \N__10318\,
            lcout => tx_shift_reg_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i8C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i10_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__10324\,
            in1 => \N__11127\,
            in2 => \N__11665\,
            in3 => \N__11052\,
            lcout => tx_shift_reg_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i8C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19_3_lut_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111011"
        )
    port map (
            in0 => \N__11716\,
            in1 => \N__12923\,
            in2 => \_gnd_net_\,
            in3 => \N__13034\,
            lcout => n5462,
            ltout => \n5462_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i6_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__10312\,
            in1 => \N__13573\,
            in2 => \N__10306\,
            in3 => \N__11076\,
            lcout => tx_shift_reg_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i7_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__10303\,
            in1 => \N__11077\,
            in2 => \N__11782\,
            in3 => \N__11126\,
            lcout => tx_shift_reg_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i251_252_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__12148\,
            in1 => \N__10288\,
            in2 => \N__10739\,
            in3 => \N__10249\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \start_tx_87_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__14318\,
            in1 => \N__10217\,
            in2 => \N__11008\,
            in3 => \N__14362\,
            lcout => \r_SM_Main_2_N_325_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i985_2_lut_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12334\,
            in2 => \_gnd_net_\,
            in3 => \N__14199\,
            lcout => rd_addr_p1_w_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i242_243_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10146\,
            in1 => \N__10724\,
            in2 => \N__10197\,
            in3 => \N__12149\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_clk_counter_i3_696__i2_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010011100"
        )
    port map (
            in0 => \N__10411\,
            in1 => \N__10382\,
            in2 => \N__10456\,
            in3 => \N__10438\,
            lcout => reset_clk_counter_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_clk_counter_i3_696__i1_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101101000100"
        )
    port map (
            in0 => \N__10437\,
            in1 => \N__10455\,
            in2 => \_gnd_net_\,
            in3 => \N__10410\,
            lcout => reset_clk_counter_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_clk_counter_i3_696__i0_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10451\,
            in2 => \_gnd_net_\,
            in3 => \N__10436\,
            lcout => reset_clk_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_all_r_81_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__10435\,
            in1 => \N__10412\,
            in2 => \N__10387\,
            in3 => \N__10368\,
            lcout => reset_all_w,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__10367\,
            in1 => \N__10381\,
            in2 => \N__10414\,
            in3 => \N__10433\,
            lcout => \reset_all_w_N_61\,
            ltout => \reset_all_w_N_61_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3898_2_lut_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__10434\,
            in1 => \_gnd_net_\,
            in2 => \N__10417\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \n2_adj_670_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_clk_counter_i3_696__i3_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101001"
        )
    port map (
            in0 => \N__10369\,
            in1 => \N__10413\,
            in2 => \N__10390\,
            in3 => \N__10386\,
            lcout => reset_clk_counter_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i1897_1_lut_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16403\,
            lcout => \RESET_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2706_2_lut_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10357\,
            in2 => \_gnd_net_\,
            in3 => \N__18932\,
            lcout => \DATA26_c_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2719_2_lut_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10801\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18936\,
            lcout => \DATA15_c_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_busy_falling_edge_83_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__10761\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10747\,
            lcout => spi_busy_falling_edge,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_busy_prev_84_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10762\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => spi_busy_prev,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.EnabledDecoder_2_i4_2_lut_3_lut_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__11249\,
            in1 => \N__12251\,
            in2 => \_gnd_net_\,
            in3 => \N__11956\,
            lcout => \tx_fifo.lscc_fifo_inst.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_write_cmd_85_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10630\,
            in2 => \_gnd_net_\,
            in3 => \N__11250\,
            lcout => fifo_write_cmd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.EnabledDecoder_2_i3_2_lut_3_lut_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__11248\,
            in1 => \N__12250\,
            in2 => \_gnd_net_\,
            in3 => \N__11955\,
            lcout => \tx_fifo.lscc_fifo_inst.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Clock_Count_700__i0_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10501\,
            in2 => \_gnd_net_\,
            in3 => \N__10489\,
            lcout => \pc_tx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \pc_tx.n4865\,
            clk => \N__19358\,
            ce => \N__16094\,
            sr => \N__10861\
        );

    \pc_tx.r_Clock_Count_700__i1_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10486\,
            in2 => \_gnd_net_\,
            in3 => \N__10474\,
            lcout => \pc_tx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \pc_tx.n4865\,
            carryout => \pc_tx.n4866\,
            clk => \N__19358\,
            ce => \N__16094\,
            sr => \N__10861\
        );

    \pc_tx.r_Clock_Count_700__i2_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10471\,
            in2 => \_gnd_net_\,
            in3 => \N__10459\,
            lcout => \pc_tx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \pc_tx.n4866\,
            carryout => \pc_tx.n4867\,
            clk => \N__19358\,
            ce => \N__16094\,
            sr => \N__10861\
        );

    \pc_tx.r_Clock_Count_700__i3_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10966\,
            in2 => \_gnd_net_\,
            in3 => \N__10954\,
            lcout => \pc_tx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \pc_tx.n4867\,
            carryout => \pc_tx.n4868\,
            clk => \N__19358\,
            ce => \N__16094\,
            sr => \N__10861\
        );

    \pc_tx.r_Clock_Count_700__i4_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10951\,
            in2 => \_gnd_net_\,
            in3 => \N__10939\,
            lcout => \pc_tx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \pc_tx.n4868\,
            carryout => \pc_tx.n4869\,
            clk => \N__19358\,
            ce => \N__16094\,
            sr => \N__10861\
        );

    \pc_tx.r_Clock_Count_700__i5_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10936\,
            in2 => \_gnd_net_\,
            in3 => \N__10924\,
            lcout => \pc_tx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \pc_tx.n4869\,
            carryout => \pc_tx.n4870\,
            clk => \N__19358\,
            ce => \N__16094\,
            sr => \N__10861\
        );

    \pc_tx.r_Clock_Count_700__i6_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10921\,
            in2 => \_gnd_net_\,
            in3 => \N__10909\,
            lcout => \pc_tx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \pc_tx.n4870\,
            carryout => \pc_tx.n4871\,
            clk => \N__19358\,
            ce => \N__16094\,
            sr => \N__10861\
        );

    \pc_tx.r_Clock_Count_700__i7_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10906\,
            in2 => \_gnd_net_\,
            in3 => \N__10894\,
            lcout => \pc_tx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \pc_tx.n4871\,
            carryout => \pc_tx.n4872\,
            clk => \N__19358\,
            ce => \N__16094\,
            sr => \N__10861\
        );

    \pc_tx.r_Clock_Count_700__i8_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10891\,
            in2 => \_gnd_net_\,
            in3 => \N__10879\,
            lcout => \pc_tx.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \pc_tx.n4873\,
            clk => \N__19354\,
            ce => \N__16095\,
            sr => \N__10857\
        );

    \pc_tx.r_Clock_Count_700__i9_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10873\,
            in2 => \_gnd_net_\,
            in3 => \N__10876\,
            lcout => \pc_tx.r_Clock_Count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19354\,
            ce => \N__16095\,
            sr => \N__10857\
        );

    \spi0.tx_shift_reg_i15_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__11137\,
            in1 => \N__11749\,
            in2 => \N__11082\,
            in3 => \N__11191\,
            lcout => \DEBUG_9_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i15C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i12_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__11218\,
            in1 => \N__11064\,
            in2 => \N__11452\,
            in3 => \N__11134\,
            lcout => tx_shift_reg_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i15C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_en_i_I_0_2_lut_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11236\,
            in2 => \_gnd_net_\,
            in3 => \N__12260\,
            lcout => wr_fifo_en_w,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i2_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__11014\,
            in1 => \N__11075\,
            in2 => \N__13804\,
            in3 => \N__11139\,
            lcout => tx_shift_reg_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i15C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i13_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__11135\,
            in1 => \N__11203\,
            in2 => \N__11081\,
            in3 => \N__11620\,
            lcout => tx_shift_reg_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i15C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i14_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__11197\,
            in1 => \N__11068\,
            in2 => \N__13597\,
            in3 => \N__11136\,
            lcout => tx_shift_reg_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i15C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i1_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__11138\,
            in1 => \N__12823\,
            in2 => \N__11083\,
            in3 => \N__11590\,
            lcout => tx_shift_reg_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i15C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_read_cmd_86_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11007\,
            in2 => \_gnd_net_\,
            in3 => \N__14319\,
            lcout => fifo_read_cmd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4497_4_lut_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111110"
        )
    port map (
            in0 => \N__14351\,
            in1 => \N__11346\,
            in2 => \N__12121\,
            in3 => \N__12336\,
            lcout => OPEN,
            ltout => \n5454_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_adj_79_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10969\,
            in3 => \N__11247\,
            lcout => OPEN,
            ltout => \n15_adj_673_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.full_r_84_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__11385\,
            in1 => \N__11635\,
            in2 => \N__11368\,
            in3 => \N__11365\,
            lcout => is_tx_fifo_full_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r__i2_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__16479\,
            in1 => \N__12204\,
            in2 => \N__11320\,
            in3 => \N__11359\,
            lcout => \tx_fifo.lscc_fifo_inst.rd_addr_r_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i1_4_lut_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001000"
        )
    port map (
            in0 => \N__11358\,
            in1 => \N__11347\,
            in2 => \N__12412\,
            in3 => \N__11644\,
            lcout => n4892,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i992_3_lut_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__12335\,
            in1 => \N__11357\,
            in2 => \_gnd_net_\,
            in3 => \N__14246\,
            lcout => rd_addr_p1_w_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_addr_r_1__I_0_i1_2_lut_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11936\,
            in2 => \_gnd_net_\,
            in3 => \N__14208\,
            lcout => n1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_en_i_I_0_2_lut_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__14352\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14298\,
            lcout => \tx_fifo.lscc_fifo_inst.rd_fifo_en_w\,
            ltout => \tx_fifo.lscc_fifo_inst.rd_fifo_en_w_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r__i1_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__16415\,
            in1 => \N__12349\,
            in2 => \N__11293\,
            in3 => \N__12220\,
            lcout => rd_addr_r_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i7_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__11849\,
            in1 => \N__11265\,
            in2 => \N__11290\,
            in3 => \N__16414\,
            lcout => fifo_temp_output_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_addr_r__i0_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000111001110"
        )
    port map (
            in0 => \N__12268\,
            in1 => \N__16427\,
            in2 => \N__11254\,
            in3 => \N__11951\,
            lcout => wr_addr_r_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19346\,
            ce => 'H',
            sr => \N__16558\
        );

    \bluejay_data_inst.i2705_2_lut_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18933\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11569\,
            lcout => \DATA27_c_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2712_2_lut_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11533\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18934\,
            lcout => \DATA20_c_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2723_2_lut_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11488\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18935\,
            lcout => \DATA13_c_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_SM_Main_i0_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__13317\,
            in1 => \N__11425\,
            in2 => \_gnd_net_\,
            in3 => \N__12664\,
            lcout => \r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19379\,
            ce => 'H',
            sr => \N__13400\
        );

    \pc_rx.r_SM_Main_i1_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001011110010"
        )
    port map (
            in0 => \N__13449\,
            in1 => \N__11431\,
            in2 => \N__13339\,
            in3 => \N__13501\,
            lcout => \r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19379\,
            ce => 'H',
            sr => \N__13400\
        );

    \tx_addr_byte_r_i0_i4_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12468\,
            in1 => \N__11442\,
            in2 => \_gnd_net_\,
            in3 => \N__15054\,
            lcout => tx_addr_byte_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i4493_2_lut_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11812\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18039\,
            lcout => \pc_rx.n5450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__18038\,
            in1 => \N__13446\,
            in2 => \_gnd_net_\,
            in3 => \N__11811\,
            lcout => \pc_rx.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i1_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11586\,
            in1 => \N__11412\,
            in2 => \_gnd_net_\,
            in3 => \N__15087\,
            lcout => tx_addr_byte_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19366\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i0_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__12489\,
            in1 => \N__18073\,
            in2 => \N__13617\,
            in3 => \N__13832\,
            lcout => pc_data_rx_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19366\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i7_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12655\,
            in1 => \N__11765\,
            in2 => \_gnd_net_\,
            in3 => \N__15090\,
            lcout => tx_data_byte_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19366\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i5_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15088\,
            in1 => \N__12431\,
            in2 => \_gnd_net_\,
            in3 => \N__11613\,
            lcout => tx_addr_byte_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19366\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i1_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__18074\,
            in1 => \N__12490\,
            in2 => \N__11602\,
            in3 => \N__12643\,
            lcout => pc_data_rx_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19366\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i1_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15089\,
            in1 => \N__11601\,
            in2 => \_gnd_net_\,
            in3 => \N__11585\,
            lcout => tx_data_byte_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19366\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_2_lut_3_lut_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__12705\,
            in1 => \N__12771\,
            in2 => \_gnd_net_\,
            in3 => \N__12750\,
            lcout => \pc_rx.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i4662_4_lut_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101010101"
        )
    port map (
            in0 => \N__13402\,
            in1 => \N__13338\,
            in2 => \N__11791\,
            in3 => \N__13460\,
            lcout => \pc_rx.n2566\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i4495_2_lut_3_lut_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__13459\,
            in1 => \N__18053\,
            in2 => \_gnd_net_\,
            in3 => \N__11805\,
            lcout => OPEN,
            ltout => \pc_rx.n5452_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_4_lut_adj_29_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010100000001"
        )
    port map (
            in0 => \N__13401\,
            in1 => \N__13337\,
            in2 => \N__11572\,
            in3 => \N__13497\,
            lcout => \pc_rx.n2705\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i4520_2_lut_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12725\,
            in2 => \_gnd_net_\,
            in3 => \N__13644\,
            lcout => OPEN,
            ltout => \pc_rx.n5478_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i4530_4_lut_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13166\,
            in1 => \N__13142\,
            in2 => \N__11824\,
            in3 => \N__13662\,
            lcout => OPEN,
            ltout => \pc_rx.n5488_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i4_4_lut_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__13118\,
            in1 => \N__11821\,
            in2 => \N__11815\,
            in3 => \N__13680\,
            lcout => \pc_rx.r_SM_Main_2_N_252_0\,
            ltout => \pc_rx.r_SM_Main_2_N_252_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2_2_lut_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__18054\,
            in1 => \_gnd_net_\,
            in2 => \N__11794\,
            in3 => \_gnd_net_\,
            lcout => \pc_rx.n6_adj_635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i7_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11772\,
            in1 => \N__15086\,
            in2 => \_gnd_net_\,
            in3 => \N__11748\,
            lcout => tx_addr_byte_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19359\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_1_lut_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11735\,
            lcout => n989,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i2_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11655\,
            in1 => \N__15091\,
            in2 => \_gnd_net_\,
            in3 => \N__13800\,
            lcout => tx_addr_byte_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i970_3_lut_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__12015\,
            in1 => \N__12233\,
            in2 => \_gnd_net_\,
            in3 => \N__11952\,
            lcout => wr_addr_p1_w_2,
            ltout => \wr_addr_p1_w_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_addr_r__i2_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__12234\,
            in1 => \N__11633\,
            in2 => \N__11638\,
            in3 => \N__16507\,
            lcout => wr_addr_r_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_addr_r__i1_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__11634\,
            in1 => \N__12057\,
            in2 => \N__16557\,
            in3 => \N__11954\,
            lcout => wr_addr_r_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_addr_p1_w_1__I_0_i2_2_lut_3_lut_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__11953\,
            in1 => \N__12014\,
            in2 => \_gnd_net_\,
            in3 => \N__12328\,
            lcout => \tx_fifo.lscc_fifo_inst.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_66_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__12337\,
            in1 => \N__14221\,
            in2 => \N__12090\,
            in3 => \N__11944\,
            lcout => OPEN,
            ltout => \n32_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14299\,
            in2 => \N__12271\,
            in3 => \N__12267\,
            lcout => n24_adj_674,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4516_4_lut_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__12235\,
            in1 => \N__12219\,
            in2 => \N__12205\,
            in3 => \N__12034\,
            lcout => OPEN,
            ltout => \n5474_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.empty_r_85_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__11908\,
            in1 => \N__16493\,
            in2 => \N__11965\,
            in3 => \N__11962\,
            lcout => is_fifo_empty_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_78_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000000000"
        )
    port map (
            in0 => \N__11945\,
            in1 => \N__14300\,
            in2 => \N__14247\,
            in3 => \N__14353\,
            lcout => n4_adj_675,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i1_2_lut_3_lut_4_lut_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__14301\,
            in1 => \N__16434\,
            in2 => \N__11833\,
            in3 => \N__14363\,
            lcout => n2545,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_fifo_en_prev_r_86_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__14302\,
            in1 => \N__16435\,
            in2 => \_gnd_net_\,
            in3 => \N__14364\,
            lcout => \tx_fifo.lscc_fifo_inst.rd_fifo_en_prev_r\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2708_2_lut_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12595\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18886\,
            lcout => \DATA24_c_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2731_2_lut_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18870\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12559\,
            lcout => \DATA5_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2730_2_lut_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12526\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18871\,
            lcout => \DATA6_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.equal_145_i4_2_lut_LC_13_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14019\,
            in2 => \_gnd_net_\,
            in3 => \N__13938\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i4_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__15052\,
            in1 => \_gnd_net_\,
            in2 => \N__12679\,
            in3 => \N__12467\,
            lcout => tx_data_byte_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2_3_lut_LC_13_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__14023\,
            in1 => \N__13942\,
            in2 => \_gnd_net_\,
            in3 => \N__12607\,
            lcout => n2468,
            ltout => \n2468_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i5_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__18041\,
            in1 => \N__12447\,
            in2 => \N__12451\,
            in3 => \N__13981\,
            lcout => pc_data_rx_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i3_LC_13_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12630\,
            in1 => \N__15051\,
            in2 => \_gnd_net_\,
            in3 => \N__13763\,
            lcout => tx_data_byte_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i5_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__15053\,
            in1 => \_gnd_net_\,
            in2 => \N__12435\,
            in3 => \N__12448\,
            lcout => tx_data_byte_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_SM_Main_i2_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__13448\,
            in1 => \N__13399\,
            in2 => \N__13354\,
            in3 => \N__13496\,
            lcout => \r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i4_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__18040\,
            in1 => \N__13980\,
            in2 => \N__12678\,
            in3 => \N__12685\,
            lcout => pc_data_rx_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_LC_13_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101101010101"
        )
    port map (
            in0 => \N__13447\,
            in1 => \N__13516\,
            in2 => \_gnd_net_\,
            in3 => \N__13495\,
            lcout => \pc_rx.n3803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_2_lut_adj_27_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__13976\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12606\,
            lcout => n2475,
            ltout => \n2475_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i7_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__13548\,
            in1 => \N__12654\,
            in2 => \N__12658\,
            in3 => \N__18072\,
            lcout => pc_data_rx_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i3_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__18071\,
            in1 => \N__13848\,
            in2 => \N__12631\,
            in3 => \N__12642\,
            lcout => pc_data_rx_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_2_lut_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12770\,
            in2 => \_gnd_net_\,
            in3 => \N__12749\,
            lcout => OPEN,
            ltout => \pc_rx.n2465_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2_4_lut_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__12704\,
            in1 => \N__12726\,
            in2 => \N__12616\,
            in3 => \N__13627\,
            lcout => OPEN,
            ltout => \pc_rx.n4887_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2904_4_lut_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__13120\,
            in1 => \N__13167\,
            in2 => \N__12613\,
            in3 => \N__13147\,
            lcout => \r_SM_Main_2_N_246_2\,
            ltout => \r_SM_Main_2_N_246_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2_3_lut_4_lut_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__13389\,
            in1 => \N__13461\,
            in2 => \N__12610\,
            in3 => \N__13336\,
            lcout => \pc_rx.n2429\,
            ltout => \pc_rx.n2429_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_2_lut_adj_28_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12781\,
            in3 => \N__13975\,
            lcout => n2471,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Clock_Count_698__i0_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13645\,
            in2 => \_gnd_net_\,
            in3 => \N__12778\,
            lcout => \pc_rx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \bfn_13_6_0_\,
            carryout => \pc_rx.n4807\,
            clk => \N__19367\,
            ce => \N__13095\,
            sr => \N__13077\
        );

    \pc_rx.r_Clock_Count_698__i1_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13681\,
            in2 => \_gnd_net_\,
            in3 => \N__12775\,
            lcout => \pc_rx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \pc_rx.n4807\,
            carryout => \pc_rx.n4808\,
            clk => \N__19367\,
            ce => \N__13095\,
            sr => \N__13077\
        );

    \pc_rx.r_Clock_Count_698__i2_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12772\,
            in2 => \_gnd_net_\,
            in3 => \N__12754\,
            lcout => \pc_rx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \pc_rx.n4808\,
            carryout => \pc_rx.n4809\,
            clk => \N__19367\,
            ce => \N__13095\,
            sr => \N__13077\
        );

    \pc_rx.r_Clock_Count_698__i3_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12751\,
            in2 => \_gnd_net_\,
            in3 => \N__12733\,
            lcout => \pc_rx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \pc_rx.n4809\,
            carryout => \pc_rx.n4810\,
            clk => \N__19367\,
            ce => \N__13095\,
            sr => \N__13077\
        );

    \pc_rx.r_Clock_Count_698__i4_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13663\,
            in2 => \_gnd_net_\,
            in3 => \N__12730\,
            lcout => \pc_rx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \pc_rx.n4810\,
            carryout => \pc_rx.n4811\,
            clk => \N__19367\,
            ce => \N__13095\,
            sr => \N__13077\
        );

    \pc_rx.r_Clock_Count_698__i5_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12727\,
            in2 => \_gnd_net_\,
            in3 => \N__12709\,
            lcout => \pc_rx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \pc_rx.n4811\,
            carryout => \pc_rx.n4812\,
            clk => \N__19367\,
            ce => \N__13095\,
            sr => \N__13077\
        );

    \pc_rx.r_Clock_Count_698__i6_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12706\,
            in2 => \_gnd_net_\,
            in3 => \N__12688\,
            lcout => \pc_rx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \pc_rx.n4812\,
            carryout => \pc_rx.n4813\,
            clk => \N__19367\,
            ce => \N__13095\,
            sr => \N__13077\
        );

    \pc_rx.r_Clock_Count_698__i7_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13168\,
            in2 => \_gnd_net_\,
            in3 => \N__13150\,
            lcout => \pc_rx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \pc_rx.n4813\,
            carryout => \pc_rx.n4814\,
            clk => \N__19367\,
            ce => \N__13095\,
            sr => \N__13077\
        );

    \pc_rx.r_Clock_Count_698__i8_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13146\,
            in2 => \_gnd_net_\,
            in3 => \N__13126\,
            lcout => \pc_rx.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \pc_rx.n4815\,
            clk => \N__19363\,
            ce => \N__13099\,
            sr => \N__13078\
        );

    \pc_rx.r_Clock_Count_698__i9_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13119\,
            in2 => \_gnd_net_\,
            in3 => \N__13123\,
            lcout => \pc_rx.r_Clock_Count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19363\,
            ce => \N__13099\,
            sr => \N__13078\
        );

    \spi0.tx_shift_reg_i0_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__13729\,
            in1 => \N__13052\,
            in2 => \_gnd_net_\,
            in3 => \N__12968\,
            lcout => tx_shift_reg_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i0C_net\,
            ce => 'H',
            sr => \N__12811\
        );

    \bluejay_data_inst.i2682_4_lut_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__18424\,
            in1 => \N__13858\,
            in2 => \N__17493\,
            in3 => \N__13267\,
            lcout => \bluejay_data_inst.n1675\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.mux_506_i4_3_lut_4_lut_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__17487\,
            in1 => \N__17149\,
            in2 => \N__18267\,
            in3 => \N__13260\,
            lcout => OPEN,
            ltout => \bluejay_data_inst.n1040_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.mux_694_i4_3_lut_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__17226\,
            in1 => \_gnd_net_\,
            in2 => \N__12796\,
            in3 => \N__17907\,
            lcout => \bluejay_data_inst.state_timeout_counter_7_N_122_3\,
            ltout => \bluejay_data_inst.state_timeout_counter_7_N_122_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i3391_4_lut_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__18255\,
            in1 => \N__17842\,
            in2 => \N__12793\,
            in3 => \N__17227\,
            lcout => OPEN,
            ltout => \bluejay_data_inst.n8_adj_656_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i1_4_lut_adj_58_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__18426\,
            in1 => \N__18592\,
            in2 => \N__12790\,
            in3 => \N__12787\,
            lcout => \bluejay_data_inst.n4_adj_648\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.mux_506_i3_3_lut_4_lut_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__17486\,
            in1 => \N__17164\,
            in2 => \N__18266\,
            in3 => \N__13259\,
            lcout => OPEN,
            ltout => \bluejay_data_inst.n1041_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.mux_694_i3_3_lut_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17906\,
            in2 => \N__13276\,
            in3 => \N__17725\,
            lcout => \bluejay_data_inst.state_timeout_counter_7_N_122_2\,
            ltout => \bluejay_data_inst.state_timeout_counter_7_N_122_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i3378_4_lut_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__13687\,
            in1 => \N__18591\,
            in2 => \N__13273\,
            in3 => \N__18425\,
            lcout => \bluejay_data_inst.n4260\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i7_4_lut_adj_55_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__14804\,
            in1 => \N__14648\,
            in2 => \N__14971\,
            in3 => \N__14510\,
            lcout => OPEN,
            ltout => \bluejay_data_inst.n18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i9_4_lut_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14939\,
            in1 => \N__14777\,
            in2 => \N__13270\,
            in3 => \N__14678\,
            lcout => \bluejay_data_inst.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i4629_2_lut_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__13261\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18264\,
            lcout => \bluejay_data_inst.n5524\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2735_2_lut_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18812\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13246\,
            lcout => \DATA1_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2711_2_lut_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18872\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13210\,
            lcout => \DATA21_c_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2_2_lut_3_lut_LC_14_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__14009\,
            in1 => \N__13974\,
            in2 => \_gnd_net_\,
            in3 => \N__13927\,
            lcout => n3753,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i4614_2_lut_3_lut_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__13462\,
            in1 => \N__13514\,
            in2 => \_gnd_net_\,
            in3 => \N__13492\,
            lcout => OPEN,
            ltout => \pc_rx.n5522_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_4_lut_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000110001"
        )
    port map (
            in0 => \N__13340\,
            in1 => \N__13392\,
            in2 => \N__13522\,
            in3 => \N__13463\,
            lcout => \pc_rx.n2676\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2781_2_lut_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13935\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14017\,
            lcout => n3672,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i4690_3_lut_4_lut_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100011"
        )
    port map (
            in0 => \N__13493\,
            in1 => \N__13390\,
            in2 => \N__13352\,
            in3 => \N__13464\,
            lcout => n5482,
            ltout => \n5482_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Bit_Index_i0_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000101100"
        )
    port map (
            in0 => \N__13348\,
            in1 => \N__13977\,
            in2 => \N__13519\,
            in3 => \N__13515\,
            lcout => \r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i13_3_lut_4_lut_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000001111"
        )
    port map (
            in0 => \N__13494\,
            in1 => \N__13391\,
            in2 => \N__13353\,
            in3 => \N__13465\,
            lcout => OPEN,
            ltout => \n2502_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_DV_52_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__13393\,
            in1 => \N__13879\,
            in2 => \N__13357\,
            in3 => \N__13347\,
            lcout => debug_led3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.equal_142_i4_2_lut_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14016\,
            in2 => \_gnd_net_\,
            in3 => \N__13934\,
            lcout => n4_adj_666,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.state_timeout_counter_i0_i5_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__15405\,
            in1 => \N__14570\,
            in2 => \_gnd_net_\,
            in3 => \N__15259\,
            lcout => \usb_to_bluejay_if_inst.state_timeout_counter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19381\,
            ce => \N__15213\,
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.state_timeout_counter_i0_i3_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__15408\,
            in1 => \N__14569\,
            in2 => \_gnd_net_\,
            in3 => \N__15298\,
            lcout => \usb_to_bluejay_if_inst.state_timeout_counter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19381\,
            ce => \N__15213\,
            sr => \_gnd_net_\
        );

    \pc_rx.i1_3_lut_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__13679\,
            in1 => \N__13661\,
            in2 => \_gnd_net_\,
            in3 => \N__13643\,
            lcout => \pc_rx.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i1_2_lut_adj_25_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15680\,
            in2 => \_gnd_net_\,
            in3 => \N__15757\,
            lcout => \usb_to_bluejay_if_inst.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i0_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13621\,
            in1 => \N__15059\,
            in2 => \_gnd_net_\,
            in3 => \N__13721\,
            lcout => tx_data_byte_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i1_2_lut_adj_16_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15404\,
            in2 => \_gnd_net_\,
            in3 => \N__15758\,
            lcout => OPEN,
            ltout => \usb_to_bluejay_if_inst.n5438_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.data_in_fifo_prev_44_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__15681\,
            in1 => \N__19560\,
            in2 => \N__13600\,
            in3 => \N__14399\,
            lcout => data_in_fifo_prev,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i6_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__15058\,
            in1 => \_gnd_net_\,
            in2 => \N__13569\,
            in3 => \N__13584\,
            lcout => tx_addr_byte_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i6_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13533\,
            in1 => \N__13562\,
            in2 => \_gnd_net_\,
            in3 => \N__15060\,
            lcout => tx_data_byte_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i6_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__13549\,
            in1 => \N__18075\,
            in2 => \N__13534\,
            in3 => \N__13833\,
            lcout => pc_data_rx_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i2_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__18079\,
            in1 => \N__13852\,
            in2 => \N__13816\,
            in3 => \N__13837\,
            lcout => pc_data_rx_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i2_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15085\,
            in1 => \N__13815\,
            in2 => \_gnd_net_\,
            in3 => \N__13793\,
            lcout => tx_data_byte_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000010"
        )
    port map (
            in0 => \N__14401\,
            in1 => \N__15691\,
            in2 => \N__19556\,
            in3 => \N__15769\,
            lcout => n10_adj_671,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i3_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15084\,
            in1 => \N__13770\,
            in2 => \_gnd_net_\,
            in3 => \N__13740\,
            lcout => tx_addr_byte_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.state__i2_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001011001100"
        )
    port map (
            in0 => \N__15407\,
            in1 => \N__15770\,
            in2 => \N__15710\,
            in3 => \N__14530\,
            lcout => state_2_adj_657,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i0_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15083\,
            in1 => \N__13698\,
            in2 => \_gnd_net_\,
            in3 => \N__13722\,
            lcout => tx_addr_byte_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i4608_2_lut_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__16828\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17721\,
            lcout => \bluejay_data_inst.n5531\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.v_counter_i10_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14941\,
            in1 => \N__14920\,
            in2 => \_gnd_net_\,
            in3 => \N__16651\,
            lcout => \bluejay_data_inst.v_counter_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19360\,
            ce => 'H',
            sr => \N__16573\
        );

    \bluejay_data_inst.v_counter_i1_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16652\,
            in1 => \N__14815\,
            in2 => \_gnd_net_\,
            in3 => \N__14833\,
            lcout => \bluejay_data_inst.v_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19360\,
            ce => 'H',
            sr => \N__16573\
        );

    \bluejay_data_inst.v_counter_i7_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14653\,
            in1 => \N__14632\,
            in2 => \_gnd_net_\,
            in3 => \N__16658\,
            lcout => \bluejay_data_inst.v_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19360\,
            ce => 'H',
            sr => \N__16573\
        );

    \bluejay_data_inst.v_counter_i2_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__14788\,
            in1 => \_gnd_net_\,
            in2 => \N__16663\,
            in3 => \N__14806\,
            lcout => \bluejay_data_inst.v_counter_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19360\,
            ce => 'H',
            sr => \N__16573\
        );

    \bluejay_data_inst.v_counter_i9_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14950\,
            in1 => \N__16659\,
            in2 => \_gnd_net_\,
            in3 => \N__14970\,
            lcout => \bluejay_data_inst.v_counter_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19360\,
            ce => 'H',
            sr => \N__16573\
        );

    \bluejay_data_inst.v_counter_i0_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16650\,
            in1 => \N__14485\,
            in2 => \_gnd_net_\,
            in3 => \N__14512\,
            lcout => \bluejay_data_inst.v_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19360\,
            ce => 'H',
            sr => \N__16573\
        );

    \bluejay_data_inst.v_counter_i6_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14680\,
            in1 => \N__14662\,
            in2 => \_gnd_net_\,
            in3 => \N__16657\,
            lcout => \bluejay_data_inst.v_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19360\,
            ce => 'H',
            sr => \N__16573\
        );

    \bluejay_data_inst.v_counter_i3_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16656\,
            in1 => \N__14761\,
            in2 => \_gnd_net_\,
            in3 => \N__14779\,
            lcout => \bluejay_data_inst.v_counter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19360\,
            ce => 'H',
            sr => \N__16573\
        );

    \bluejay_data_inst.i8_4_lut_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14618\,
            in1 => \N__14831\,
            in2 => \N__14712\,
            in3 => \N__14744\,
            lcout => \bluejay_data_inst.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.v_counter_i4_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__14745\,
            in1 => \_gnd_net_\,
            in2 => \N__14731\,
            in3 => \N__16645\,
            lcout => \bluejay_data_inst.v_counter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19351\,
            ce => 'H',
            sr => \N__16567\
        );

    \bluejay_data_inst.v_counter_i8_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14622\,
            in1 => \N__14602\,
            in2 => \_gnd_net_\,
            in3 => \N__16649\,
            lcout => \bluejay_data_inst.v_counter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19351\,
            ce => 'H',
            sr => \N__16567\
        );

    \bluejay_data_inst.v_counter_i5_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__14708\,
            in1 => \_gnd_net_\,
            in2 => \N__16662\,
            in3 => \N__14692\,
            lcout => \bluejay_data_inst.v_counter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19351\,
            ce => 'H',
            sr => \N__16567\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r__i0_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000110101110"
        )
    port map (
            in0 => \N__16572\,
            in1 => \N__14368\,
            in2 => \N__14320\,
            in3 => \N__14198\,
            lcout => rd_addr_r_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19351\,
            ce => 'H',
            sr => \N__16567\
        );

    \bluejay_data_inst.i2726_2_lut_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14149\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18811\,
            lcout => \DATA10_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2727_2_lut_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14110\,
            in2 => \_gnd_net_\,
            in3 => \N__18882\,
            lcout => \DATA9_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2718_2_lut_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14068\,
            in2 => \_gnd_net_\,
            in3 => \N__18931\,
            lcout => \DATA16_c_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Bit_Index_i2_LC_15_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__13937\,
            in1 => \N__14018\,
            in2 => \_gnd_net_\,
            in3 => \N__13979\,
            lcout => \pc_rx.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19393\,
            ce => \N__13900\,
            sr => \N__13894\
        );

    \pc_rx.r_Bit_Index_i1_LC_15_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13978\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13936\,
            lcout => \pc_rx.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19393\,
            ce => \N__13900\,
            sr => \N__13894\
        );

    \uart_rx_complete_prev_89_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13878\,
            lcout => uart_rx_complete_prev,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_start_transfer_r_90_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14989\,
            in2 => \_gnd_net_\,
            in3 => \N__15021\,
            lcout => spi_start_transfer_r,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_complete_rising_edge_88_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13877\,
            in2 => \_gnd_net_\,
            in3 => \N__13864\,
            lcout => uart_rx_complete_rising_edge,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.start_transfer_edge_73_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__14418\,
            in1 => \N__14407\,
            in2 => \N__14476\,
            in3 => \N__14436\,
            lcout => start_transfer_edge,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i5_4_lut_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15309\,
            in1 => \N__15270\,
            in2 => \N__15229\,
            in3 => \N__15246\,
            lcout => \usb_to_bluejay_if_inst.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i103_2_lut_3_lut_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__15400\,
            in1 => \N__15707\,
            in2 => \_gnd_net_\,
            in3 => \N__15781\,
            lcout => \usb_to_bluejay_if_inst.n81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i2_3_lut_4_lut_adj_20_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__14392\,
            in1 => \N__14563\,
            in2 => \N__19566\,
            in3 => \N__15399\,
            lcout => \usb_to_bluejay_if_inst.n5400\,
            ltout => \usb_to_bluejay_if_inst.n5400_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i2_3_lut_4_lut_adj_15_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__15401\,
            in1 => \N__15708\,
            in2 => \N__14425\,
            in3 => \N__15782\,
            lcout => \usb_to_bluejay_if_inst.n2527\,
            ltout => \usb_to_bluejay_if_inst.n2527_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i1_4_lut_4_lut_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__15783\,
            in1 => \N__15709\,
            in2 => \N__14422\,
            in3 => \N__15402\,
            lcout => \usb_to_bluejay_if_inst.n4120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.start_transfer_prev_74_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14419\,
            lcout => start_transfer_prev,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i3253_3_lut_4_lut_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110000"
        )
    port map (
            in0 => \N__15811\,
            in1 => \N__19561\,
            in2 => \N__14400\,
            in3 => \N__15390\,
            lcout => OPEN,
            ltout => \usb_to_bluejay_if_inst.n4136_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i1_3_lut_4_lut_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__15598\,
            in1 => \N__15615\,
            in2 => \N__14371\,
            in3 => \N__14572\,
            lcout => \usb_to_bluejay_if_inst.n2492\,
            ltout => \usb_to_bluejay_if_inst.n2492_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i2_4_lut_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__15755\,
            in1 => \N__15702\,
            in2 => \N__14593\,
            in3 => \N__15392\,
            lcout => \usb_to_bluejay_if_inst.n4963\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.state__i0_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__15393\,
            in1 => \N__15756\,
            in2 => \N__15712\,
            in3 => \N__15812\,
            lcout => state_0_adj_658,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19382\,
            ce => \N__14590\,
            sr => \N__14581\
        );

    \usb_to_bluejay_if_inst.i1_2_lut_3_lut_adj_23_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__15753\,
            in1 => \N__15701\,
            in2 => \_gnd_net_\,
            in3 => \N__15388\,
            lcout => \usb_to_bluejay_if_inst.state_timeout_counter_7__N_178\,
            ltout => \usb_to_bluejay_if_inst.state_timeout_counter_7__N_178_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i2_3_lut_4_lut_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__15389\,
            in1 => \N__14571\,
            in2 => \N__14542\,
            in3 => \N__15810\,
            lcout => OPEN,
            ltout => \usb_to_bluejay_if_inst.n2562_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i1_4_lut_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__15616\,
            in1 => \N__14539\,
            in2 => \N__14533\,
            in3 => \N__15597\,
            lcout => \usb_to_bluejay_if_inst.n2564\,
            ltout => \usb_to_bluejay_if_inst.n2564_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i1_3_lut_4_lut_adj_24_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__15391\,
            in1 => \N__15706\,
            in2 => \N__14524\,
            in3 => \N__15754\,
            lcout => \usb_to_bluejay_if_inst.n2706\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.state__i1_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__15406\,
            in1 => \N__15771\,
            in2 => \N__15711\,
            in3 => \N__15814\,
            lcout => state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19374\,
            ce => \N__15322\,
            sr => \N__14521\
        );

    \bluejay_data_inst.i2693_2_lut_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14869\,
            in2 => \N__14909\,
            in3 => \N__17494\,
            lcout => \bluejay_data_inst.n1476\,
            ltout => OPEN,
            carryin => \bfn_15_8_0_\,
            carryout => \bluejay_data_inst.n4847\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.add_692_2_lut_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14511\,
            in2 => \N__14494\,
            in3 => \N__14479\,
            lcout => \bluejay_data_inst.n1109\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4847\,
            carryout => \bluejay_data_inst.n4848\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.add_692_3_lut_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14832\,
            in2 => \N__14910\,
            in3 => \N__14809\,
            lcout => \bluejay_data_inst.n1108\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4848\,
            carryout => \bluejay_data_inst.n4849\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.add_692_4_lut_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14805\,
            in2 => \N__14895\,
            in3 => \N__14782\,
            lcout => \bluejay_data_inst.n1107\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4849\,
            carryout => \bluejay_data_inst.n4850\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.add_692_5_lut_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14778\,
            in2 => \N__14911\,
            in3 => \N__14755\,
            lcout => \bluejay_data_inst.n1106\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4850\,
            carryout => \bluejay_data_inst.n4851\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.add_692_6_lut_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14752\,
            in2 => \N__14896\,
            in3 => \N__14719\,
            lcout => \bluejay_data_inst.n1105\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4851\,
            carryout => \bluejay_data_inst.n4852\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.add_692_7_lut_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14876\,
            in2 => \N__14716\,
            in3 => \N__14683\,
            lcout => \bluejay_data_inst.n1104\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4852\,
            carryout => \bluejay_data_inst.n4853\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.add_692_8_lut_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14679\,
            in2 => \N__14897\,
            in3 => \N__14656\,
            lcout => \bluejay_data_inst.n1103\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4853\,
            carryout => \bluejay_data_inst.n4854\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.add_692_9_lut_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14649\,
            in2 => \N__14907\,
            in3 => \N__14626\,
            lcout => \bluejay_data_inst.n1102\,
            ltout => OPEN,
            carryin => \bfn_15_9_0_\,
            carryout => \bluejay_data_inst.n4855\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.add_692_10_lut_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14890\,
            in2 => \N__14623\,
            in3 => \N__14596\,
            lcout => \bluejay_data_inst.n1101\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4855\,
            carryout => \bluejay_data_inst.n4856\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.add_692_11_lut_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14969\,
            in2 => \N__14908\,
            in3 => \N__14944\,
            lcout => \bluejay_data_inst.n1100\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4856\,
            carryout => \bluejay_data_inst.n4857\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.add_692_12_lut_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14894\,
            in1 => \N__14940\,
            in2 => \_gnd_net_\,
            in3 => \N__14923\,
            lcout => \bluejay_data_inst.n1099\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i1206_2_lut_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__16642\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16524\,
            lcout => \bluejay_data_inst.n2096\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i12_3_lut_3_lut_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001000100"
        )
    port map (
            in0 => \N__18364\,
            in1 => \N__18504\,
            in2 => \_gnd_net_\,
            in3 => \N__18167\,
            lcout => \bluejay_data_inst.n1054\,
            ltout => \bluejay_data_inst.n1054_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2_2_lut_3_lut_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__18168\,
            in1 => \_gnd_net_\,
            in2 => \N__14914\,
            in3 => \N__18365\,
            lcout => \bluejay_data_inst.n1373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i680_2_lut_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17899\,
            in2 => \_gnd_net_\,
            in3 => \N__17488\,
            lcout => \bluejay_data_inst.n1432\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.state__i1_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100110000"
        )
    port map (
            in0 => \N__16644\,
            in1 => \N__15961\,
            in2 => \N__18435\,
            in3 => \N__17524\,
            lcout => \bluejay_data_inst.state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19356\,
            ce => 'H',
            sr => \N__16568\
        );

    \bluejay_data_inst.i1727_2_lut_3_lut_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__18505\,
            in1 => \N__18388\,
            in2 => \_gnd_net_\,
            in3 => \N__18181\,
            lcout => n5,
            ltout => \n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.state__i0_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__17523\,
            in1 => \N__17419\,
            in2 => \N__14836\,
            in3 => \N__15967\,
            lcout => state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19356\,
            ce => 'H',
            sr => \N__16568\
        );

    \bluejay_data_inst.i1804_4_lut_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__16829\,
            in1 => \N__16566\,
            in2 => \N__17549\,
            in3 => \N__16698\,
            lcout => \bluejay_data_inst.n2693\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.state__i2_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__15187\,
            in1 => \N__16643\,
            in2 => \N__15178\,
            in3 => \N__18506\,
            lcout => state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19356\,
            ce => 'H',
            sr => \N__16568\
        );

    \bluejay_data_inst.i2733_2_lut_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18760\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15169\,
            lcout => \DATA3_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.equal_558_i3_2_lut_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18371\,
            in2 => \_gnd_net_\,
            in3 => \N__18509\,
            lcout => n3_adj_669,
            ltout => \n3_adj_669_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_75_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111010"
        )
    port map (
            in0 => \N__16492\,
            in1 => \N__16640\,
            in2 => \N__15127\,
            in3 => \N__18200\,
            lcout => n2555,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2724_2_lut_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18759\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15124\,
            lcout => \DATA12_c_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \even_byte_flag_95_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14988\,
            in2 => \_gnd_net_\,
            in3 => \N__15022\,
            lcout => even_byte_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.state_timeout_counter_i0_i0_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15835\,
            in2 => \_gnd_net_\,
            in3 => \N__14977\,
            lcout => \usb_to_bluejay_if_inst.state_timeout_counter_0\,
            ltout => OPEN,
            carryin => \bfn_16_5_0_\,
            carryout => \usb_to_bluejay_if_inst.n4800\,
            clk => \N__19391\,
            ce => \N__15214\,
            sr => \N__15196\
        );

    \usb_to_bluejay_if_inst.state_timeout_counter_i0_i1_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15859\,
            in2 => \N__17034\,
            in3 => \N__14974\,
            lcout => \usb_to_bluejay_if_inst.state_timeout_counter_1\,
            ltout => OPEN,
            carryin => \usb_to_bluejay_if_inst.n4800\,
            carryout => \usb_to_bluejay_if_inst.n4801\,
            clk => \N__19391\,
            ce => \N__15214\,
            sr => \N__15196\
        );

    \usb_to_bluejay_if_inst.state_timeout_counter_i0_i2_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15871\,
            in2 => \N__17037\,
            in3 => \N__15316\,
            lcout => \usb_to_bluejay_if_inst.state_timeout_counter_2\,
            ltout => OPEN,
            carryin => \usb_to_bluejay_if_inst.n4801\,
            carryout => \usb_to_bluejay_if_inst.n4802\,
            clk => \N__19391\,
            ce => \N__15214\,
            sr => \N__15196\
        );

    \usb_to_bluejay_if_inst.sub_123_add_2_5_lut_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__15283\,
            in1 => \N__15313\,
            in2 => \N__17035\,
            in3 => \N__15289\,
            lcout => \usb_to_bluejay_if_inst.n82\,
            ltout => OPEN,
            carryin => \usb_to_bluejay_if_inst.n4802\,
            carryout => \usb_to_bluejay_if_inst.n4803\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.state_timeout_counter_i0_i4_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15847\,
            in2 => \N__17038\,
            in3 => \N__15286\,
            lcout => \usb_to_bluejay_if_inst.state_timeout_counter_4\,
            ltout => OPEN,
            carryin => \usb_to_bluejay_if_inst.n4803\,
            carryout => \usb_to_bluejay_if_inst.n4804\,
            clk => \N__19391\,
            ce => \N__15214\,
            sr => \N__15196\
        );

    \usb_to_bluejay_if_inst.sub_123_add_2_7_lut_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__15282\,
            in1 => \N__15274\,
            in2 => \N__17036\,
            in3 => \N__15250\,
            lcout => \usb_to_bluejay_if_inst.n83\,
            ltout => OPEN,
            carryin => \usb_to_bluejay_if_inst.n4804\,
            carryout => \usb_to_bluejay_if_inst.n4805\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.state_timeout_counter_i0_i6_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15247\,
            in2 => \N__17039\,
            in3 => \N__15235\,
            lcout => \usb_to_bluejay_if_inst.state_timeout_counter_6\,
            ltout => OPEN,
            carryin => \usb_to_bluejay_if_inst.n4805\,
            carryout => \usb_to_bluejay_if_inst.n4806\,
            clk => \N__19391\,
            ce => \N__15214\,
            sr => \N__15196\
        );

    \usb_to_bluejay_if_inst.state_timeout_counter_i0_i7_LC_16_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15228\,
            in1 => \N__16997\,
            in2 => \_gnd_net_\,
            in3 => \N__15232\,
            lcout => \usb_to_bluejay_if_inst.state_timeout_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19391\,
            ce => \N__15214\,
            sr => \N__15196\
        );

    \usb_to_bluejay_if_inst.i4631_2_lut_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15983\,
            in2 => \_gnd_net_\,
            in3 => \N__18655\,
            lcout => n5546,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.next_line_rdy_o_40_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__15685\,
            in1 => \N__15398\,
            in2 => \_gnd_net_\,
            in3 => \N__15787\,
            lcout => \DEBUG_3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i23_4_lut_4_lut_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001010100"
        )
    port map (
            in0 => \N__15786\,
            in1 => \N__15684\,
            in2 => \N__15409\,
            in3 => \N__15813\,
            lcout => n16_adj_672,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i4_2_lut_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15870\,
            in2 => \_gnd_net_\,
            in3 => \N__15858\,
            lcout => OPEN,
            ltout => \usb_to_bluejay_if_inst.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i7_4_lut_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__15846\,
            in1 => \N__15834\,
            in2 => \N__15823\,
            in3 => \N__15820\,
            lcout => n11,
            ltout => \n11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i104_3_lut_4_lut_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001010"
        )
    port map (
            in0 => \N__15682\,
            in1 => \N__15394\,
            in2 => \N__15790\,
            in3 => \N__15784\,
            lcout => OPEN,
            ltout => \usb_to_bluejay_if_inst.n82_adj_628_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i2_3_lut_4_lut_adj_18_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110001"
        )
    port map (
            in0 => \N__15785\,
            in1 => \N__15683\,
            in2 => \N__15619\,
            in3 => \N__15614\,
            lcout => \usb_to_bluejay_if_inst.n2561\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_SM_Main_i2_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__15589\,
            in1 => \N__16147\,
            in2 => \N__15544\,
            in3 => \N__15463\,
            lcout => \r_SM_Main_2_adj_659\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.h_counter__i3_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__17550\,
            in1 => \N__16858\,
            in2 => \N__18265\,
            in3 => \N__17780\,
            lcout => \bluejay_data_inst.h_counter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19383\,
            ce => \N__16716\,
            sr => \N__16579\
        );

    \bluejay_data_inst.h_counter__i5_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__18245\,
            in1 => \N__17551\,
            in2 => \N__17782\,
            in3 => \N__16765\,
            lcout => \bluejay_data_inst.h_counter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19383\,
            ce => \N__16716\,
            sr => \N__16579\
        );

    \i1_3_lut_adj_70_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__15424\,
            in1 => \N__15415\,
            in2 => \_gnd_net_\,
            in3 => \N__15403\,
            lcout => n5122,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i6_4_lut_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16776\,
            in1 => \N__16752\,
            in2 => \N__16735\,
            in3 => \N__16845\,
            lcout => OPEN,
            ltout => \bluejay_data_inst.n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i7_4_lut_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__16033\,
            in1 => \N__16051\,
            in2 => \N__15904\,
            in3 => \N__15886\,
            lcout => \bluejay_data_inst.valid_o_N_155\,
            ltout => \bluejay_data_inst.valid_o_N_155_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.get_next_word_cmd_82_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__17522\,
            in1 => \N__15901\,
            in2 => \N__15889\,
            in3 => \N__18419\,
            lcout => get_next_word_cmd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19375\,
            ce => 'H',
            sr => \N__17503\
        );

    \bluejay_data_inst.i2_2_lut_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__16869\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16884\,
            lcout => \bluejay_data_inst.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i1_2_lut_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16815\,
            in2 => \_gnd_net_\,
            in3 => \N__18418\,
            lcout => \bluejay_data_inst.n31\,
            ltout => \bluejay_data_inst.n31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i3371_4_lut_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__18601\,
            in1 => \N__17316\,
            in2 => \N__15880\,
            in3 => \N__15954\,
            lcout => OPEN,
            ltout => \bluejay_data_inst.n4253_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i3374_4_lut_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__15955\,
            in1 => \N__17772\,
            in2 => \N__15877\,
            in3 => \N__18244\,
            lcout => \bluejay_data_inst.n4_adj_652\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.mux_506_i6_3_lut_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__18179\,
            in1 => \N__17131\,
            in2 => \_gnd_net_\,
            in3 => \N__17480\,
            lcout => OPEN,
            ltout => \bluejay_data_inst.n1038_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.mux_694_i6_3_lut_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__17901\,
            in1 => \_gnd_net_\,
            in2 => \N__15874\,
            in3 => \N__17409\,
            lcout => \bluejay_data_inst.state_timeout_counter_7_N_122_5\,
            ltout => \bluejay_data_inst.state_timeout_counter_7_N_122_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i3384_4_lut_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__17410\,
            in1 => \N__16012\,
            in2 => \N__16006\,
            in3 => \N__18508\,
            lcout => \bluejay_data_inst.n4266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i3401_4_lut_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110100"
        )
    port map (
            in0 => \N__16817\,
            in1 => \N__18372\,
            in2 => \N__15996\,
            in3 => \N__18180\,
            lcout => \bluejay_data_inst.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2_3_lut_adj_51_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__16641\,
            in1 => \N__17902\,
            in2 => \_gnd_net_\,
            in3 => \N__17481\,
            lcout => \bluejay_data_inst.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i1_2_lut_adj_35_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16816\,
            in2 => \_gnd_net_\,
            in3 => \N__18507\,
            lcout => \bluejay_data_inst.n34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i3370_3_lut_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17900\,
            in1 => \N__16672\,
            in2 => \_gnd_net_\,
            in3 => \N__17315\,
            lcout => \bluejay_data_inst.n4252\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.state_timeout_counter_i3_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__18546\,
            in1 => \N__18413\,
            in2 => \_gnd_net_\,
            in3 => \N__17212\,
            lcout => \bluejay_data_inst.state_timeout_counter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19361\,
            ce => 'H',
            sr => \N__15946\
        );

    \bluejay_data_inst.i32_4_lut_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__16830\,
            in1 => \N__18544\,
            in2 => \N__15927\,
            in3 => \N__18379\,
            lcout => OPEN,
            ltout => \bluejay_data_inst.n3627_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.valid_o_79_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110110000"
        )
    port map (
            in0 => \N__15923\,
            in1 => \N__16661\,
            in2 => \N__15934\,
            in3 => \N__18206\,
            lcout => \VALID_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19369\,
            ce => 'H',
            sr => \N__16577\
        );

    \bluejay_data_inst.i32_4_lut_adj_48_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011110000"
        )
    port map (
            in0 => \N__16831\,
            in1 => \N__18545\,
            in2 => \N__18810\,
            in3 => \N__18380\,
            lcout => OPEN,
            ltout => \bluejay_data_inst.n3631_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.data_output_active_cmd_84_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110110000"
        )
    port map (
            in0 => \N__18758\,
            in1 => \N__16660\,
            in2 => \N__16582\,
            in3 => \N__18205\,
            lcout => \bluejay_data_inst.data_output_active_cmd\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19369\,
            ce => 'H',
            sr => \N__16577\
        );

    \bluejay_data_inst.i3387_4_lut_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__16318\,
            in1 => \N__18204\,
            in2 => \N__17773\,
            in3 => \N__16309\,
            lcout => \bluejay_data_inst.n4_adj_637\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.state_timeout_counter_i1_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__18587\,
            in1 => \N__18423\,
            in2 => \_gnd_net_\,
            in3 => \N__17310\,
            lcout => \bluejay_data_inst.state_timeout_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19376\,
            ce => 'H',
            sr => \N__16300\
        );

    \bluejay_data_inst.i2672_2_lut_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18828\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16291\,
            lcout => \DATA0_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2710_2_lut_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16239\,
            in2 => \_gnd_net_\,
            in3 => \N__18919\,
            lcout => \DEBUG_5_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i1_1_lut_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16140\,
            lcout => \pc_tx.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.h_counter__i0_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16050\,
            in2 => \_gnd_net_\,
            in3 => \N__16036\,
            lcout => \bluejay_data_inst.h_counter_0\,
            ltout => OPEN,
            carryin => \bfn_17_7_0_\,
            carryout => \bluejay_data_inst.n4858\,
            clk => \N__19387\,
            ce => \N__16717\,
            sr => \N__16687\
        );

    \bluejay_data_inst.h_counter__i1_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16032\,
            in2 => \N__17040\,
            in3 => \N__16015\,
            lcout => \bluejay_data_inst.h_counter_1\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4858\,
            carryout => \bluejay_data_inst.n4859\,
            clk => \N__19387\,
            ce => \N__16717\,
            sr => \N__16687\
        );

    \bluejay_data_inst.h_counter__i2_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17001\,
            in2 => \N__16891\,
            in3 => \N__16873\,
            lcout => \bluejay_data_inst.h_counter_2\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4859\,
            carryout => \bluejay_data_inst.n4860\,
            clk => \N__19387\,
            ce => \N__16717\,
            sr => \N__16687\
        );

    \bluejay_data_inst.sub_117_add_2_5_lut_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16821\,
            in1 => \N__16870\,
            in2 => \N__17041\,
            in3 => \N__16852\,
            lcout => \bluejay_data_inst.n5547\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4860\,
            carryout => \bluejay_data_inst.n4861\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.h_counter__i4_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17002\,
            in2 => \N__16849\,
            in3 => \N__16834\,
            lcout => \bluejay_data_inst.h_counter_4\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4861\,
            carryout => \bluejay_data_inst.n4862\,
            clk => \N__19387\,
            ce => \N__16717\,
            sr => \N__16687\
        );

    \bluejay_data_inst.sub_117_add_2_7_lut_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16822\,
            in1 => \N__16777\,
            in2 => \N__17042\,
            in3 => \N__16759\,
            lcout => \bluejay_data_inst.n5548\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4862\,
            carryout => \bluejay_data_inst.n4863\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.h_counter__i6_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17003\,
            in2 => \N__16756\,
            in3 => \N__16741\,
            lcout => \bluejay_data_inst.h_counter_6\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4863\,
            carryout => \bluejay_data_inst.n4864\,
            clk => \N__19387\,
            ce => \N__16717\,
            sr => \N__16687\
        );

    \bluejay_data_inst.h_counter__i7_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17004\,
            in1 => \N__16731\,
            in2 => \_gnd_net_\,
            in3 => \N__16738\,
            lcout => \bluejay_data_inst.h_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19387\,
            ce => \N__16717\,
            sr => \N__16687\
        );

    \bluejay_data_inst.sub_119_add_2_2_lut_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17475\,
            in1 => \N__17671\,
            in2 => \_gnd_net_\,
            in3 => \N__16675\,
            lcout => \bluejay_data_inst.n5521\,
            ltout => OPEN,
            carryin => \bfn_17_8_0_\,
            carryout => \bluejay_data_inst.n4816\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.sub_119_add_2_3_lut_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17476\,
            in1 => \N__17317\,
            in2 => \N__17055\,
            in3 => \N__16666\,
            lcout => \bluejay_data_inst.n5527\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4816\,
            carryout => \bluejay_data_inst.n4817\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.sub_119_add_2_4_lut_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17714\,
            in2 => \N__17061\,
            in3 => \N__17152\,
            lcout => \bluejay_data_inst.n51\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4817\,
            carryout => \bluejay_data_inst.n4818\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.sub_119_add_2_5_lut_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17225\,
            in2 => \N__17056\,
            in3 => \N__17137\,
            lcout => \bluejay_data_inst.n50\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4818\,
            carryout => \bluejay_data_inst.n4819\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.sub_119_add_2_6_lut_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17248\,
            in2 => \N__17062\,
            in3 => \N__17134\,
            lcout => \bluejay_data_inst.n49\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4819\,
            carryout => \bluejay_data_inst.n4820\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.sub_119_add_2_7_lut_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17407\,
            in2 => \N__17057\,
            in3 => \N__17125\,
            lcout => \bluejay_data_inst.n48\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4820\,
            carryout => \bluejay_data_inst.n4821\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.sub_119_add_2_8_lut_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17474\,
            in1 => \N__17967\,
            in2 => \N__17063\,
            in3 => \N__17122\,
            lcout => \bluejay_data_inst.n5545\,
            ltout => OPEN,
            carryin => \bluejay_data_inst.n4821\,
            carryout => \bluejay_data_inst.n4822\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.sub_119_add_2_9_lut_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__17030\,
            in1 => \N__17587\,
            in2 => \N__17492\,
            in3 => \N__16906\,
            lcout => \bluejay_data_inst.n5544\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.mux_694_i5_3_lut_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17249\,
            in1 => \N__17903\,
            in2 => \_gnd_net_\,
            in3 => \N__17266\,
            lcout => \bluejay_data_inst.state_timeout_counter_7_N_122_4\,
            ltout => \bluejay_data_inst.state_timeout_counter_7_N_122_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i3395_4_lut_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__17823\,
            in1 => \N__18257\,
            in2 => \N__16903\,
            in3 => \N__17250\,
            lcout => OPEN,
            ltout => \bluejay_data_inst.n8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i1_4_lut_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__16900\,
            in1 => \N__18593\,
            in2 => \N__16894\,
            in3 => \N__18429\,
            lcout => \bluejay_data_inst.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2_2_lut_adj_52_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17311\,
            in2 => \_gnd_net_\,
            in3 => \N__17704\,
            lcout => OPEN,
            ltout => \bluejay_data_inst.n10_adj_654_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i7_4_lut_adj_54_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__17408\,
            in1 => \N__17672\,
            in2 => \N__17278\,
            in3 => \N__17191\,
            lcout => \bluejay_data_inst.n1394\,
            ltout => \bluejay_data_inst.n1394_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.mux_506_i5_3_lut_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101111"
        )
    port map (
            in0 => \N__17275\,
            in1 => \_gnd_net_\,
            in2 => \N__17269\,
            in3 => \N__18256\,
            lcout => \bluejay_data_inst.n1039\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.state_timeout_counter_i4_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__17251\,
            in1 => \N__18594\,
            in2 => \_gnd_net_\,
            in3 => \N__18430\,
            lcout => \bluejay_data_inst.state_timeout_counter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19377\,
            ce => 'H',
            sr => \N__17260\
        );

    \bluejay_data_inst.i6_4_lut_adj_53_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17247\,
            in1 => \N__17580\,
            in2 => \N__17971\,
            in3 => \N__17224\,
            lcout => \bluejay_data_inst.n14_adj_655\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.mux_694_i8_3_lut_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17916\,
            in1 => \N__17185\,
            in2 => \_gnd_net_\,
            in3 => \N__17584\,
            lcout => \bluejay_data_inst.state_timeout_counter_7_N_122_7\,
            ltout => \bluejay_data_inst.state_timeout_counter_7_N_122_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i21_4_lut_adj_31_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__17585\,
            in1 => \N__17841\,
            in2 => \N__17176\,
            in3 => \N__18242\,
            lcout => OPEN,
            ltout => \bluejay_data_inst.n8_adj_640_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i1_4_lut_adj_32_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__18578\,
            in1 => \N__17173\,
            in2 => \N__17167\,
            in3 => \N__18390\,
            lcout => \bluejay_data_inst.n4_adj_641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.state_timeout_counter_i7_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__17586\,
            in1 => \N__18579\,
            in2 => \_gnd_net_\,
            in3 => \N__18414\,
            lcout => \bluejay_data_inst.state_timeout_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19364\,
            ce => 'H',
            sr => \N__17560\
        );

    \bluejay_data_inst.i2_2_lut_3_lut_adj_50_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__18575\,
            in1 => \N__18389\,
            in2 => \_gnd_net_\,
            in3 => \N__18231\,
            lcout => \bluejay_data_inst.n5_adj_653\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2713_2_lut_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18576\,
            in2 => \_gnd_net_\,
            in3 => \N__18243\,
            lcout => \bluejay_data_inst.n3602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i1_2_lut_3_lut_adj_22_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__18577\,
            in1 => \N__18656\,
            in2 => \_gnd_net_\,
            in3 => \N__18233\,
            lcout => n15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.mux_532_i1_3_lut_3_lut_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001100110"
        )
    port map (
            in0 => \N__18232\,
            in1 => \N__17917\,
            in2 => \_gnd_net_\,
            in3 => \N__17482\,
            lcout => \bluejay_data_inst.n1133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.state_timeout_counter_i5_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__18603\,
            in1 => \N__18434\,
            in2 => \_gnd_net_\,
            in3 => \N__17398\,
            lcout => \bluejay_data_inst.state_timeout_counter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19378\,
            ce => 'H',
            sr => \N__17371\
        );

    \bluejay_data_inst.i2732_2_lut_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18866\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17359\,
            lcout => \DATA4_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.state_timeout_counter_i6_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__18602\,
            in1 => \N__18432\,
            in2 => \_gnd_net_\,
            in3 => \N__17970\,
            lcout => \bluejay_data_inst.state_timeout_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19388\,
            ce => 'H',
            sr => \N__17929\
        );

    \bluejay_data_inst.mux_694_i7_3_lut_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17905\,
            in1 => \N__17323\,
            in2 => \_gnd_net_\,
            in3 => \N__17968\,
            lcout => \bluejay_data_inst.state_timeout_counter_7_N_122_6\,
            ltout => \bluejay_data_inst.state_timeout_counter_7_N_122_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i21_4_lut_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__17969\,
            in1 => \N__17836\,
            in2 => \N__17941\,
            in3 => \N__18258\,
            lcout => OPEN,
            ltout => \bluejay_data_inst.n8_adj_638_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i1_4_lut_adj_30_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__18427\,
            in1 => \N__17938\,
            in2 => \N__17932\,
            in3 => \N__18595\,
            lcout => \bluejay_data_inst.n4_adj_639\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.mux_694_i1_3_lut_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17904\,
            in1 => \N__17848\,
            in2 => \_gnd_net_\,
            in3 => \N__17673\,
            lcout => \bluejay_data_inst.state_timeout_counter_7_N_122_0\,
            ltout => \bluejay_data_inst.state_timeout_counter_7_N_122_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i21_4_lut_adj_36_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__17674\,
            in1 => \N__17837\,
            in2 => \N__17803\,
            in3 => \N__18262\,
            lcout => OPEN,
            ltout => \bluejay_data_inst.n8_adj_645_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i1_4_lut_adj_62_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__18596\,
            in1 => \N__18428\,
            in2 => \N__17800\,
            in3 => \N__17797\,
            lcout => \bluejay_data_inst.n4_adj_636\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i3381_4_lut_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__18263\,
            in1 => \N__17791\,
            in2 => \N__17781\,
            in3 => \N__17734\,
            lcout => \bluejay_data_inst.n4_adj_650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.state_timeout_counter_i2_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__18580\,
            in1 => \N__18431\,
            in2 => \_gnd_net_\,
            in3 => \N__17713\,
            lcout => \bluejay_data_inst.state_timeout_counter_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19370\,
            ce => 'H',
            sr => \N__17683\
        );

    \bluejay_data_inst.state_timeout_counter_i0_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__18433\,
            in1 => \N__18600\,
            in2 => \_gnd_net_\,
            in3 => \N__17659\,
            lcout => \bluejay_data_inst.state_timeout_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19392\,
            ce => 'H',
            sr => \N__17641\
        );

    \bluejay_data_inst.i2729_2_lut_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18914\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17629\,
            lcout => \DATA7_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2717_2_lut_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19009\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18915\,
            lcout => \DATA17_c_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.i2734_2_lut_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18954\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18700\,
            lcout => \DATA2_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.i3309_1_lut_2_lut_LC_19_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__18663\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19567\,
            lcout => \DEBUG_8_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bluejay_data_inst.update_o_80_LC_19_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18604\,
            in1 => \N__18436\,
            in2 => \_gnd_net_\,
            in3 => \N__18268\,
            lcout => \UPDATE_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19389\,
            ce => 'H',
            sr => \N__18091\
        );

    \pc_rx.r_Rx_Data_50_LC_20_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19417\,
            lcout => \r_Rx_Data\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19399\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i0_LC_23_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17998\,
            in2 => \_gnd_net_\,
            in3 => \N__17992\,
            lcout => n25_adj_662,
            ltout => OPEN,
            carryin => \bfn_23_5_0_\,
            carryout => n4823,
            clk => \N__19402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i1_LC_23_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17989\,
            in2 => \_gnd_net_\,
            in3 => \N__17983\,
            lcout => n24,
            ltout => OPEN,
            carryin => n4823,
            carryout => n4824,
            clk => \N__19402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i2_LC_23_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17980\,
            in2 => \_gnd_net_\,
            in3 => \N__17974\,
            lcout => n23,
            ltout => OPEN,
            carryin => n4824,
            carryout => n4825,
            clk => \N__19402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i3_LC_23_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19081\,
            in2 => \_gnd_net_\,
            in3 => \N__19075\,
            lcout => n22,
            ltout => OPEN,
            carryin => n4825,
            carryout => n4826,
            clk => \N__19402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i4_LC_23_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19072\,
            in2 => \_gnd_net_\,
            in3 => \N__19066\,
            lcout => n21,
            ltout => OPEN,
            carryin => n4826,
            carryout => n4827,
            clk => \N__19402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i5_LC_23_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19063\,
            in2 => \_gnd_net_\,
            in3 => \N__19057\,
            lcout => n20,
            ltout => OPEN,
            carryin => n4827,
            carryout => n4828,
            clk => \N__19402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i6_LC_23_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19054\,
            in2 => \_gnd_net_\,
            in3 => \N__19048\,
            lcout => n19,
            ltout => OPEN,
            carryin => n4828,
            carryout => n4829,
            clk => \N__19402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i7_LC_23_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19045\,
            in2 => \_gnd_net_\,
            in3 => \N__19039\,
            lcout => n18,
            ltout => OPEN,
            carryin => n4829,
            carryout => n4830,
            clk => \N__19402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i8_LC_23_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19036\,
            in2 => \_gnd_net_\,
            in3 => \N__19030\,
            lcout => n17,
            ltout => OPEN,
            carryin => \bfn_23_6_0_\,
            carryout => n4831,
            clk => \N__19401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i9_LC_23_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19027\,
            in2 => \_gnd_net_\,
            in3 => \N__19021\,
            lcout => n16,
            ltout => OPEN,
            carryin => n4831,
            carryout => n4832,
            clk => \N__19401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i10_LC_23_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19018\,
            in2 => \_gnd_net_\,
            in3 => \N__19012\,
            lcout => n15_adj_663,
            ltout => OPEN,
            carryin => n4832,
            carryout => n4833,
            clk => \N__19401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i11_LC_23_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19162\,
            in2 => \_gnd_net_\,
            in3 => \N__19156\,
            lcout => n14,
            ltout => OPEN,
            carryin => n4833,
            carryout => n4834,
            clk => \N__19401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i12_LC_23_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19153\,
            in2 => \_gnd_net_\,
            in3 => \N__19147\,
            lcout => n13,
            ltout => OPEN,
            carryin => n4834,
            carryout => n4835,
            clk => \N__19401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i13_LC_23_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19144\,
            in2 => \_gnd_net_\,
            in3 => \N__19138\,
            lcout => n12,
            ltout => OPEN,
            carryin => n4835,
            carryout => n4836,
            clk => \N__19401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i14_LC_23_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19135\,
            in2 => \_gnd_net_\,
            in3 => \N__19129\,
            lcout => n11_adj_661,
            ltout => OPEN,
            carryin => n4836,
            carryout => n4837,
            clk => \N__19401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i15_LC_23_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19126\,
            in2 => \_gnd_net_\,
            in3 => \N__19120\,
            lcout => n10,
            ltout => OPEN,
            carryin => n4837,
            carryout => n4838,
            clk => \N__19401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i16_LC_23_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19117\,
            in2 => \_gnd_net_\,
            in3 => \N__19111\,
            lcout => n9,
            ltout => OPEN,
            carryin => \bfn_23_7_0_\,
            carryout => n4839,
            clk => \N__19400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i17_LC_23_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19108\,
            in2 => \_gnd_net_\,
            in3 => \N__19102\,
            lcout => n8,
            ltout => OPEN,
            carryin => n4839,
            carryout => n4840,
            clk => \N__19400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i18_LC_23_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19099\,
            in2 => \_gnd_net_\,
            in3 => \N__19093\,
            lcout => n7,
            ltout => OPEN,
            carryin => n4840,
            carryout => n4841,
            clk => \N__19400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i19_LC_23_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19090\,
            in2 => \_gnd_net_\,
            in3 => \N__19084\,
            lcout => n6,
            ltout => OPEN,
            carryin => n4841,
            carryout => n4842,
            clk => \N__19400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i20_LC_23_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19630\,
            in2 => \_gnd_net_\,
            in3 => \N__19624\,
            lcout => n5_adj_665,
            ltout => OPEN,
            carryin => n4842,
            carryout => n4843,
            clk => \N__19400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i21_LC_23_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19621\,
            in2 => \_gnd_net_\,
            in3 => \N__19615\,
            lcout => n4_adj_664,
            ltout => OPEN,
            carryin => n4843,
            carryout => n4844,
            clk => \N__19400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i22_LC_23_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19612\,
            in2 => \_gnd_net_\,
            in3 => \N__19606\,
            lcout => n3,
            ltout => OPEN,
            carryin => n4844,
            carryout => n4845,
            clk => \N__19400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i23_LC_23_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19603\,
            in2 => \_gnd_net_\,
            in3 => \N__19597\,
            lcout => n2,
            ltout => OPEN,
            carryin => n4845,
            carryout => n4846,
            clk => \N__19400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_695_867__i24_LC_23_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19578\,
            in2 => \_gnd_net_\,
            in3 => \N__19594\,
            lcout => \DEBUG_0_c_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \usb_to_bluejay_if_inst.fifo_empty_i_I_0_1_lut_LC_23_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19565\,
            lcout => \DEBUG_1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_SLM_CLK_c_THRU_LUT4_0_LC_23_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19408\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_SLM_CLK_c_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Data_R_49_LC_24_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19432\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pc_rx.r_Rx_Data_R\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19403\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

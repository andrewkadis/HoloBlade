// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Thu Feb 27 21:49:18 2020
//
// Verilog Description of module top
//

module top (ICE_SYSCLK, DCD, DSR, DTR, CTS, RST, UART_RX, UART_TX, 
            SEN, SCK, SOUT, SDAT, UPDATE, RESET, SLM_CLK, INVERT, 
            SYNC, VALID, DATA31, DATA0, DATA30, DATA29, DATA1, 
            DATA28, DATA27, DATA2, DATA26, DATA25, DATA3, DATA24, 
            DATA23, DATA4, DATA22, DATA21, DATA5, DATA20, DATA19, 
            DATA6, DATA18, DATA17, DATA7, DATA16, DATA15, DATA8, 
            DATA14, DATA13, DATA12, DATA11, DATA9, DATA10, FT_OE, 
            FT_RD, FT_WR, FT_SIWU, FR_RXF, FT_TXE, FIFO_BE3, FIFO_BE2, 
            FIFO_BE1, FIFO_BE0, FIFO_D31, FIFO_D30, FIFO_D29, FIFO_D28, 
            FIFO_D27, FIFO_CLK, FIFO_D26, FIFO_D25, FIFO_D24, FIFO_D23, 
            FIFO_D22, FIFO_D21, FIFO_D20, FIFO_D19, FIFO_D18, FIFO_D17, 
            FIFO_D16, FIFO_D15, FIFO_D14, FIFO_D13, FIFO_D12, FIFO_D11, 
            FIFO_D10, FIFO_D9, FIFO_D8, FIFO_D7, FIFO_D6, FIFO_D5, 
            FIFO_D4, FIFO_D3, FIFO_D2, FIFO_D1, FIFO_D0, DEBUG_0, 
            DEBUG_1, DEBUG_2, DEBUG_3, DEBUG_5, DEBUG_6, DEBUG_8, 
            DEBUG_9, ICE_CLK, ICE_CDONE, ICE_CREST) /* synthesis syn_module_defined=1 */ ;   // src/top.v(5[8:11])
    input ICE_SYSCLK;   // src/top.v(8[11:21])
    output DCD;   // src/top.v(11[12:15])
    output DSR;   // src/top.v(12[12:15])
    output DTR;   // src/top.v(13[12:15])
    output CTS;   // src/top.v(14[12:15])
    output RST;   // src/top.v(15[12:15])
    input UART_RX;   // src/top.v(16[12:19])
    output UART_TX;   // src/top.v(17[12:19])
    output SEN;   // src/top.v(20[12:15])
    output SCK;   // src/top.v(21[12:15])
    input SOUT;   // src/top.v(22[12:16])
    output SDAT;   // src/top.v(23[12:16])
    output UPDATE;   // src/top.v(27[12:18])
    output RESET;   // src/top.v(28[12:17])
    output SLM_CLK;   // src/top.v(29[12:19])
    output INVERT;   // src/top.v(30[12:18])
    output SYNC;   // src/top.v(31[12:16])
    output VALID;   // src/top.v(32[12:17])
    output DATA31;   // src/top.v(34[12:18])
    output DATA0;   // src/top.v(35[12:17])
    output DATA30;   // src/top.v(36[12:18])
    output DATA29;   // src/top.v(37[12:18])
    output DATA1;   // src/top.v(38[12:17])
    output DATA28;   // src/top.v(39[12:18])
    output DATA27;   // src/top.v(40[12:18])
    output DATA2;   // src/top.v(41[12:17])
    output DATA26;   // src/top.v(42[12:18])
    output DATA25;   // src/top.v(43[12:18])
    output DATA3;   // src/top.v(44[12:17])
    output DATA24;   // src/top.v(45[12:18])
    output DATA23;   // src/top.v(46[12:18])
    output DATA4;   // src/top.v(47[12:17])
    output DATA22;   // src/top.v(48[12:18])
    output DATA21;   // src/top.v(49[12:18])
    output DATA5;   // src/top.v(50[12:17])
    output DATA20;   // src/top.v(51[12:18])
    output DATA19;   // src/top.v(52[12:18])
    output DATA6;   // src/top.v(53[12:17])
    output DATA18;   // src/top.v(54[12:18])
    output DATA17;   // src/top.v(55[12:18])
    output DATA7;   // src/top.v(56[12:17])
    output DATA16;   // src/top.v(57[12:18])
    output DATA15;   // src/top.v(58[12:18])
    output DATA8;   // src/top.v(59[12:17])
    output DATA14;   // src/top.v(60[12:18])
    output DATA13;   // src/top.v(61[12:18])
    output DATA12;   // src/top.v(62[12:18])
    output DATA11;   // src/top.v(63[12:18])
    output DATA9;   // src/top.v(64[12:17])
    output DATA10;   // src/top.v(65[12:18])
    output FT_OE;   // src/top.v(69[12:17])
    output FT_RD;   // src/top.v(70[12:17])
    output FT_WR;   // src/top.v(71[12:17])
    output FT_SIWU;   // src/top.v(72[12:19])
    input FR_RXF;   // src/top.v(73[12:18])
    input FT_TXE;   // src/top.v(74[12:18])
    output FIFO_BE3;   // src/top.v(75[12:20])
    output FIFO_BE2;   // src/top.v(76[12:20])
    output FIFO_BE1;   // src/top.v(77[12:20])
    output FIFO_BE0;   // src/top.v(78[12:20])
    output FIFO_D31;   // src/top.v(79[12:20])
    output FIFO_D30;   // src/top.v(80[12:20])
    output FIFO_D29;   // src/top.v(81[12:20])
    output FIFO_D28;   // src/top.v(82[12:20])
    output FIFO_D27;   // src/top.v(83[12:20])
    input FIFO_CLK;   // src/top.v(84[12:20])
    output FIFO_D26;   // src/top.v(85[12:20])
    output FIFO_D25;   // src/top.v(86[12:20])
    output FIFO_D24;   // src/top.v(87[12:20])
    output FIFO_D23;   // src/top.v(88[12:20])
    output FIFO_D22;   // src/top.v(89[12:20])
    output FIFO_D21;   // src/top.v(90[12:20])
    output FIFO_D20;   // src/top.v(91[12:20])
    output FIFO_D19;   // src/top.v(92[12:20])
    output FIFO_D18;   // src/top.v(93[12:20])
    output FIFO_D17;   // src/top.v(94[12:20])
    output FIFO_D16;   // src/top.v(95[12:20])
    output FIFO_D15;   // src/top.v(97[12:20])
    output FIFO_D14;   // src/top.v(98[12:20])
    output FIFO_D13;   // src/top.v(99[12:20])
    output FIFO_D12;   // src/top.v(100[12:20])
    output FIFO_D11;   // src/top.v(101[12:20])
    output FIFO_D10;   // src/top.v(102[12:20])
    output FIFO_D9;   // src/top.v(103[12:19])
    output FIFO_D8;   // src/top.v(104[12:19])
    output FIFO_D7;   // src/top.v(105[12:19])
    output FIFO_D6;   // src/top.v(106[12:19])
    output FIFO_D5;   // src/top.v(107[12:19])
    output FIFO_D4;   // src/top.v(108[12:19])
    output FIFO_D3;   // src/top.v(109[12:19])
    output FIFO_D2;   // src/top.v(110[12:19])
    output FIFO_D1;   // src/top.v(111[12:19])
    input FIFO_D0;   // src/top.v(112[12:19])
    output DEBUG_0;   // src/top.v(115[12:19])
    output DEBUG_1;   // src/top.v(116[12:19])
    output DEBUG_2;   // src/top.v(117[12:19])
    output DEBUG_3;   // src/top.v(118[12:19])
    output DEBUG_5;   // src/top.v(119[12:19])
    output DEBUG_6;   // src/top.v(120[12:19])
    output DEBUG_8;   // src/top.v(121[12:19])
    output DEBUG_9;   // src/top.v(122[12:19])
    output ICE_CLK;   // src/top.v(125[12:19])
    output ICE_CDONE;   // src/top.v(126[12:21])
    output ICE_CREST;   // src/top.v(127[12:21])
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    
    wire GND_net, VCC_net, ICE_SYSCLK_c, UART_RX_c, UART_TX_c, SEN_c, 
        DEBUG_6_c, DEBUG_5_c_c, SDAT_c, RESET_c, FT_OE_c, FT_RD_c, 
        DEBUG_9_c_c, DEBUG_8_c_c, DEBUG_0_c_24, DEBUG_1_c, DEBUG_2_c, 
        n1965, reset_all_w;
    wire [3:0]reset_clk_counter;   // src/top.v(233[10:27])
    wire [7:0]pc_data_rx;   // src/top.v(373[11:21])
    
    wire tx_uart_active_flag, spi_busy;
    wire [7:0]tx_addr_byte;   // src/top.v(485[11:23])
    wire [7:0]tx_data_byte;   // src/top.v(487[11:23])
    wire [7:0]rx_buf_byte;   // src/top.v(494[11:22])
    
    wire is_tx_fifo_full_flag, fifo_write_cmd, spi_busy_falling_edge, 
        spi_busy_prev, fifo_read_cmd, is_fifo_empty_flag;
    wire [31:0]fifo_temp_output;   // src/top.v(577[12:28])
    
    wire even_byte_flag, uart_rx_complete_rising_edge, uart_rx_complete_prev, 
        n1963, n1636, reset_all_w_N_61, n1962, n1961, r_Rx_Data, 
        start_tx_N_71, pll_clk_unbuf, n24, \mem_LUT.mem_3_7 , \mem_LUT.mem_3_6 , 
        \mem_LUT.mem_3_5 , \mem_LUT.mem_3_4 , \mem_LUT.mem_3_3 , \mem_LUT.mem_3_2 , 
        \mem_LUT.mem_3_1 , \mem_LUT.mem_3_0 ;
    wire [2:0]r_Bit_Index;   // src/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // src/uart_rx.v(36[17:26])
    
    wire n4, n8, n4_adj_494, n2, n1819, n2968;
    wire [2:0]r_SM_Main_2__N_108;
    
    wire n3178, n2540;
    wire [2:0]r_SM_Main_adj_512;   // src/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_514;   // src/uart_tx.v(33[16:27])
    wire [7:0]r_Tx_Data;   // src/uart_tx.v(34[16:25])
    wire [2:0]r_SM_Main_2__N_187;
    wire [2:0]r_SM_Main_2__N_184;
    
    wire n8_adj_499, n2959, n3206, n3190, n2076, n23, n2073;
    wire [15:0]tx_shift_reg;   // src/spi.v(66[26:38])
    wire [15:0]rx_shift_reg;   // src/spi.v(67[26:38])
    
    wire start_transfer_edge, start_transfer_prev;
    wire [2:0]state_reg;   // src/spi.v(132[10:19])
    
    wire n2068, n2067, n1957, n1956, n2066, n2065, n2064, n2958, 
        n2062, state_next_2__N_312, n2061, n2060, n2059, n2058, 
        n2057, n2056, n2055, n2054, n2053, n2052, n2051, n2050, 
        n2049, n2048, n2047, n2046, n2045, n2044, n2043, n2042, 
        rx_shift_reg_15__N_319, n2041, n2040, n2039, n2038, n2037, 
        n2036, n2035, n2034, n2033, n2032, n2031, n2030, n2029, 
        n2025, n2957, n1747, n2956, n1795, n1954, wr_fifo_en_w, 
        rd_fifo_en_w, rd_fifo_en_prev_r, n2016;
    wire [2:0]wr_addr_r;   // src/fifo_quad_word_mod.v(65[31:40])
    wire [2:0]wr_addr_p1_w;   // src/fifo_quad_word_mod.v(67[32:44])
    wire [2:0]rd_addr_r;   // src/fifo_quad_word_mod.v(69[31:40])
    wire [2:0]rd_addr_p1_w;   // src/fifo_quad_word_mod.v(71[32:44])
    
    wire n4_adj_500, n13, n12, n11, n10, n9, n8_adj_501, n7, 
        n6, n5, n4_adj_502, n3, n2_adj_503, n2955, n2013;
    wire [31:0]\mem_LUT.data_raw_r ;   // src/fifo_quad_word_mod.v(449[42:52])
    
    wire n2954, n2953, n14, n2010, n2009, n3180, n2005, n2004, 
        n2003, n2002, n2001, n2000, n1285, n1999, n1998, n1997, 
        n1996, n1995, n1994, n2952, n1951, n1950, \mem_LUT.mem_1_7 , 
        \mem_LUT.mem_1_6 , \mem_LUT.mem_1_5 , \mem_LUT.mem_1_4 , \mem_LUT.mem_1_3 , 
        \mem_LUT.mem_1_2 , n1991, n1949, n4_adj_504, n1990, n1948, 
        n2951, n1945, n1944, n2950, n1942, n1898, \mem_LUT.mem_1_1 , 
        \mem_LUT.mem_1_0 , n2949, n1988, n2948, n122, n123, n124, 
        n2947, n1983, n883, n125, n2_adj_505, n1939, n126, n127, 
        n1982, n1938, n2946, n1981, n128, n129, n130, n2945, 
        n1978, n121, n120, n119, n118, n117, n116, n115, n114, 
        n113, n112, n111, n110, n109, n108, n107, n106, n4_adj_506, 
        n1764, n19, n2944, n5_adj_507, n2943, n17, n25, n16, 
        n22, n15, n2942, n2941, n2994, n21, n18, n2992, n1, 
        n3239, n2940, n20, n1728, n1935, n1933, n1930, n1929, 
        n1975, n1974, n1973, n1972, n1971, n1968, n2939, n25_adj_508, 
        n2938, n2990, n2961, n1754, n1750, n2960, n3118, n15_adj_509, 
        n3275, n24_adj_510, n32, n3279, n4_adj_511, n3148, n3448, 
        n3250, n3439, n3184, n3188, n3198, n3293, n3204, n3289, 
        n3212;
    
    VCC i2 (.Y(VCC_net));
    spi spi0 (.state_reg({state_reg}), .state_next_2__N_312(state_next_2__N_312), 
        .VCC_net(VCC_net), .SDAT_c(SDAT_c), .reset_all_w(reset_all_w), 
        .DEBUG_2_c(DEBUG_2_c), .start_transfer_prev(start_transfer_prev), 
        .SLM_CLK_c(SLM_CLK_c), .n3212(n3212), .\rx_shift_reg[8] (rx_shift_reg[8]), 
        .\tx_shift_reg[0] (tx_shift_reg[0]), .n3206(n3206), .\rx_shift_reg[7] (rx_shift_reg[7]), 
        .n3204(n3204), .\rx_shift_reg[6] (rx_shift_reg[6]), .n3198(n3198), 
        .\rx_shift_reg[5] (rx_shift_reg[5]), .SEN_c(SEN_c), .n3190(n3190), 
        .\rx_shift_reg[4] (rx_shift_reg[4]), .n3188(n3188), .\rx_shift_reg[3] (rx_shift_reg[3]), 
        .n3184(n3184), .\rx_shift_reg[2] (rx_shift_reg[2]), .n3180(n3180), 
        .\rx_shift_reg[1] (rx_shift_reg[1]), .n2059(n2059), .\tx_shift_reg[1] (tx_shift_reg[1]), 
        .n2057(n2057), .\tx_shift_reg[2] (tx_shift_reg[2]), .n2055(n2055), 
        .\tx_shift_reg[3] (tx_shift_reg[3]), .n2054(n2054), .\tx_shift_reg[4] (tx_shift_reg[4]), 
        .n2053(n2053), .\tx_shift_reg[5] (tx_shift_reg[5]), .n2052(n2052), 
        .\tx_shift_reg[6] (tx_shift_reg[6]), .n2043(n2043), .\tx_shift_reg[7] (tx_shift_reg[7]), 
        .n2042(n2042), .\tx_shift_reg[8] (tx_shift_reg[8]), .n2041(n2041), 
        .\tx_shift_reg[9] (tx_shift_reg[9]), .n2040(n2040), .\tx_shift_reg[10] (tx_shift_reg[10]), 
        .n2039(n2039), .\tx_shift_reg[11] (tx_shift_reg[11]), .n2038(n2038), 
        .\tx_shift_reg[12] (tx_shift_reg[12]), .n2037(n2037), .\tx_shift_reg[13] (tx_shift_reg[13]), 
        .n2036(n2036), .n2034(n2034), .rx_buf_byte({rx_buf_byte}), .n2033(n2033), 
        .n2032(n2032), .n2031(n2031), .n2030(n2030), .n3148(n3148), 
        .start_transfer_edge(start_transfer_edge), .n2029(n2029), .n2025(n2025), 
        .GND_net(GND_net), .spi_busy(spi_busy), .n1956(n1956), .n3178(n3178), 
        .\rx_shift_reg[0] (rx_shift_reg[0]), .n1728(n1728), .n5(n5_adj_507), 
        .DEBUG_6_c(DEBUG_6_c), .rx_shift_reg_15__N_319(rx_shift_reg_15__N_319), 
        .\tx_data_byte[0] (tx_data_byte[0]), .n883(n883), .n3279(n3279), 
        .\tx_addr_byte[7] (tx_addr_byte[7])) /* synthesis syn_module_defined=1 */ ;   // src/top.v(511[5] 534[2])
    SB_DFF reset_all_r_198 (.Q(reset_all_w), .C(SLM_CLK_c), .D(reset_all_w_N_61));   // src/top.v(237[8] 255[4])
    SB_DFF spi_busy_prev_203 (.Q(spi_busy_prev), .C(SLM_CLK_c), .D(spi_busy));   // src/top.v(552[8] 558[4])
    SB_DFF fifo_read_cmd_205 (.Q(fifo_read_cmd), .C(SLM_CLK_c), .D(start_tx_N_71));   // src/top.v(581[8] 599[4])
    SB_DFF uart_rx_complete_prev_208 (.Q(uart_rx_complete_prev), .C(SLM_CLK_c), 
           .D(DEBUG_1_c));   // src/top.v(739[8] 745[4])
    SB_IO RST_pad (.PACKAGE_PIN(RST), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RST_pad.PIN_TYPE = 6'b011001;
    defparam RST_pad.PULLUP = 1'b0;
    defparam RST_pad.NEG_TRIGGER = 1'b0;
    defparam RST_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB clk_gb (.GLOBAL_BUFFER_OUTPUT(SLM_CLK_c), .USER_SIGNAL_TO_GLOBAL_BUFFER(pll_clk_unbuf)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=214, LSE_RLINE=219 */ ;   // src/clock.v(30[7:96])
    SB_DFF led_counter_581_788__i0 (.Q(n25), .C(SLM_CLK_c), .D(n130));   // src/top.v(195[20:35])
    SB_IO UART_TX_pad (.PACKAGE_PIN(UART_TX), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(UART_TX_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UART_TX_pad.PIN_TYPE = 6'b011001;
    defparam UART_TX_pad.PULLUP = 1'b0;
    defparam UART_TX_pad.NEG_TRIGGER = 1'b0;
    defparam UART_TX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA31_pad (.PACKAGE_PIN(DATA31), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA31_pad.PIN_TYPE = 6'b011001;
    defparam DATA31_pad.PULLUP = 1'b0;
    defparam DATA31_pad.NEG_TRIGGER = 1'b0;
    defparam DATA31_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1695_3_lut (.I0(\mem_LUT.mem_3_4 ), .I1(rx_buf_byte[4]), .I2(n2), 
            .I3(GND_net), .O(n2048));   // src/fifo_quad_word_mod.v(448[73:76])
    defparam i1695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1612_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[3]), .I2(n4_adj_504), 
            .I3(n1754), .O(n1965));   // src/uart_rx.v(49[10] 144[8])
    defparam i1612_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1696_3_lut (.I0(\mem_LUT.mem_3_5 ), .I1(rx_buf_byte[5]), .I2(n2), 
            .I3(GND_net), .O(n2049));   // src/fifo_quad_word_mod.v(448[73:76])
    defparam i1696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1697_3_lut (.I0(\mem_LUT.mem_3_6 ), .I1(rx_buf_byte[6]), .I2(n2), 
            .I3(GND_net), .O(n2050));   // src/fifo_quad_word_mod.v(448[73:76])
    defparam i1697_3_lut.LUT_INIT = 16'hcaca;
    SB_IO VALID_pad (.PACKAGE_PIN(VALID), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam VALID_pad.PIN_TYPE = 6'b011001;
    defparam VALID_pad.PULLUP = 1'b0;
    defparam VALID_pad.NEG_TRIGGER = 1'b0;
    defparam VALID_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1698_3_lut (.I0(\mem_LUT.mem_3_7 ), .I1(rx_buf_byte[7]), .I2(n2), 
            .I3(GND_net), .O(n2051));   // src/fifo_quad_word_mod.v(448[73:76])
    defparam i1698_3_lut.LUT_INIT = 16'hcaca;
    SB_IO SYNC_pad (.PACKAGE_PIN(SYNC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SYNC_pad.PIN_TYPE = 6'b011001;
    defparam SYNC_pad.PULLUP = 1'b0;
    defparam SYNC_pad.NEG_TRIGGER = 1'b0;
    defparam SYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INVERT_pad (.PACKAGE_PIN(INVERT), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INVERT_pad.PIN_TYPE = 6'b011001;
    defparam INVERT_pad.PULLUP = 1'b0;
    defparam INVERT_pad.NEG_TRIGGER = 1'b0;
    defparam INVERT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SLM_CLK_pad (.PACKAGE_PIN(SLM_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SLM_CLK_c));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SLM_CLK_pad.PIN_TYPE = 6'b011001;
    defparam SLM_CLK_pad.PULLUP = 1'b0;
    defparam SLM_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam SLM_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFF even_byte_flag_214 (.Q(even_byte_flag), .C(SLM_CLK_c), .D(n1285));   // src/top.v(748[8] 802[4])
    SB_IO RESET_pad (.PACKAGE_PIN(RESET), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(RESET_c));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RESET_pad.PIN_TYPE = 6'b011001;
    defparam RESET_pad.PULLUP = 1'b0;
    defparam RESET_pad.NEG_TRIGGER = 1'b0;
    defparam RESET_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UPDATE_pad (.PACKAGE_PIN(UPDATE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UPDATE_pad.PIN_TYPE = 6'b011001;
    defparam UPDATE_pad.PULLUP = 1'b0;
    defparam UPDATE_pad.NEG_TRIGGER = 1'b0;
    defparam UPDATE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SDAT_pad (.PACKAGE_PIN(SDAT), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SDAT_c));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SDAT_pad.PIN_TYPE = 6'b011001;
    defparam SDAT_pad.PULLUP = 1'b0;
    defparam SDAT_pad.NEG_TRIGGER = 1'b0;
    defparam SDAT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SCK_pad (.PACKAGE_PIN(SCK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_6_c));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SCK_pad.PIN_TYPE = 6'b011001;
    defparam SCK_pad.PULLUP = 1'b0;
    defparam SCK_pad.NEG_TRIGGER = 1'b0;
    defparam SCK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SEN_pad (.PACKAGE_PIN(SEN), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SEN_c));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SEN_pad.PIN_TYPE = 6'b011001;
    defparam SEN_pad.PULLUP = 1'b0;
    defparam SEN_pad.NEG_TRIGGER = 1'b0;
    defparam SEN_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CTS_pad (.PACKAGE_PIN(CTS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CTS_pad.PIN_TYPE = 6'b011001;
    defparam CTS_pad.PULLUP = 1'b0;
    defparam CTS_pad.NEG_TRIGGER = 1'b0;
    defparam CTS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY led_counter_581_788_add_4_21 (.CI(n2956), .I0(GND_net), .I1(n6), 
            .CO(n2957));
    SB_LUT4 i1_2_lut (.I0(rx_shift_reg[5]), .I1(n3279), .I2(GND_net), 
            .I3(GND_net), .O(n3204));   // src/spi.v(299[8] 313[4])
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1699_4_lut (.I0(tx_shift_reg[5]), .I1(tx_data_byte[6]), .I2(n3279), 
            .I3(n1728), .O(n2052));   // src/spi.v(275[8] 290[4])
    defparam i1699_4_lut.LUT_INIT = 16'hce0a;
    SB_IO DTR_pad (.PACKAGE_PIN(DTR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DTR_pad.PIN_TYPE = 6'b011001;
    defparam DTR_pad.PULLUP = 1'b0;
    defparam DTR_pad.NEG_TRIGGER = 1'b0;
    defparam DTR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DSR_pad (.PACKAGE_PIN(DSR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DSR_pad.PIN_TYPE = 6'b011001;
    defparam DSR_pad.PULLUP = 1'b0;
    defparam DSR_pad.NEG_TRIGGER = 1'b0;
    defparam DSR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DCD_pad (.PACKAGE_PIN(DCD), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DCD_pad.PIN_TYPE = 6'b011001;
    defparam DCD_pad.PULLUP = 1'b0;
    defparam DCD_pad.NEG_TRIGGER = 1'b0;
    defparam DCD_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFF tx_data_byte_r_i0_i1 (.Q(tx_data_byte[1]), .C(SLM_CLK_c), .D(n2068));   // src/top.v(748[8] 802[4])
    SB_IO DATA0_pad (.PACKAGE_PIN(DATA0), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA0_pad.PIN_TYPE = 6'b011001;
    defparam DATA0_pad.PULLUP = 1'b0;
    defparam DATA0_pad.NEG_TRIGGER = 1'b0;
    defparam DATA0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1619_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[4]), .I2(n4_adj_506), 
            .I3(n1750), .O(n1972));   // src/uart_rx.v(49[10] 144[8])
    defparam i1619_4_lut.LUT_INIT = 16'hccca;
    SB_DFF tx_addr_byte_r_i0_i0 (.Q(tx_addr_byte[0]), .C(SLM_CLK_c), .D(n1961));   // src/top.v(748[8] 802[4])
    SB_DFF tx_data_byte_r_i0_i2 (.Q(tx_data_byte[2]), .C(SLM_CLK_c), .D(n2058));   // src/top.v(748[8] 802[4])
    SB_DFF reset_clk_counter_i3_582__i0 (.Q(reset_clk_counter[0]), .C(SLM_CLK_c), 
           .D(n25_adj_508));   // src/top.v(250[27:51])
    SB_DFF tx_data_byte_r_i0_i3 (.Q(tx_data_byte[3]), .C(SLM_CLK_c), .D(n2056));   // src/top.v(748[8] 802[4])
    SB_LUT4 i1620_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[5]), .I2(n4_adj_506), 
            .I3(n1754), .O(n1973));   // src/uart_rx.v(49[10] 144[8])
    defparam i1620_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1621_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[6]), .I2(r_Bit_Index[0]), 
            .I3(n1747), .O(n1974));   // src/uart_rx.v(49[10] 144[8])
    defparam i1621_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY led_counter_581_788_add_4_11 (.CI(n2946), .I0(GND_net), .I1(n16), 
            .CO(n2947));
    SB_LUT4 led_counter_581_788_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17), .I3(n2945), .O(n122)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_18 (.I0(rx_shift_reg[6]), .I1(n3279), .I2(GND_net), 
            .I3(GND_net), .O(n3206));   // src/spi.v(299[8] 313[4])
    defparam i1_2_lut_adj_18.LUT_INIT = 16'h2222;
    SB_CARRY led_counter_581_788_add_4_10 (.CI(n2945), .I0(GND_net), .I1(n17), 
            .CO(n2946));
    SB_LUT4 led_counter_581_788_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18), .I3(n2944), .O(n123)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1622_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[7]), .I2(r_Bit_Index[0]), 
            .I3(n1747), .O(n1975));   // src/uart_rx.v(49[10] 144[8])
    defparam i1622_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1629_2_lut (.I0(uart_rx_complete_rising_edge), .I1(even_byte_flag), 
            .I2(GND_net), .I3(GND_net), .O(n1982));   // src/top.v(748[8] 802[4])
    defparam i1629_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1628_4_lut_4_lut (.I0(rd_fifo_en_w), .I1(reset_all_w), .I2(rd_addr_p1_w[2]), 
            .I3(rd_addr_r[2]), .O(n1981));
    defparam i1628_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_DFF led_counter_581_788__i24 (.Q(DEBUG_0_c_24), .C(SLM_CLK_c), .D(n106));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i23 (.Q(n2_adj_503), .C(SLM_CLK_c), .D(n107));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i22 (.Q(n3), .C(SLM_CLK_c), .D(n108));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i21 (.Q(n4_adj_502), .C(SLM_CLK_c), .D(n109));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i20 (.Q(n5), .C(SLM_CLK_c), .D(n110));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i19 (.Q(n6), .C(SLM_CLK_c), .D(n111));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i18 (.Q(n7), .C(SLM_CLK_c), .D(n112));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i17 (.Q(n8_adj_501), .C(SLM_CLK_c), .D(n113));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i16 (.Q(n9), .C(SLM_CLK_c), .D(n114));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i15 (.Q(n10), .C(SLM_CLK_c), .D(n115));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i14 (.Q(n11), .C(SLM_CLK_c), .D(n116));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i13 (.Q(n12), .C(SLM_CLK_c), .D(n117));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i12 (.Q(n13), .C(SLM_CLK_c), .D(n118));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i11 (.Q(n14), .C(SLM_CLK_c), .D(n119));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i10 (.Q(n15), .C(SLM_CLK_c), .D(n120));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i9 (.Q(n16), .C(SLM_CLK_c), .D(n121));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i8 (.Q(n17), .C(SLM_CLK_c), .D(n122));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i7 (.Q(n18), .C(SLM_CLK_c), .D(n123));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i6 (.Q(n19), .C(SLM_CLK_c), .D(n124));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i5 (.Q(n20), .C(SLM_CLK_c), .D(n125));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i4 (.Q(n21), .C(SLM_CLK_c), .D(n126));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i3 (.Q(n22), .C(SLM_CLK_c), .D(n127));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i2 (.Q(n23), .C(SLM_CLK_c), .D(n128));   // src/top.v(195[20:35])
    SB_DFF led_counter_581_788__i1 (.Q(n24), .C(SLM_CLK_c), .D(n129));   // src/top.v(195[20:35])
    SB_DFF FT_RD_r_201 (.Q(FT_RD_c), .C(FIFO_CLK_c), .D(FT_OE_c));   // src/top.v(289[8] 303[6])
    SB_LUT4 i1625_4_lut_4_lut (.I0(rd_fifo_en_w), .I1(reset_all_w), .I2(rd_addr_r[0]), 
            .I3(rd_addr_r[1]), .O(n1978));
    defparam i1625_4_lut_4_lut.LUT_INIT = 16'h1320;
    SB_LUT4 i1700_4_lut (.I0(tx_shift_reg[4]), .I1(tx_data_byte[5]), .I2(n3279), 
            .I3(n1728), .O(n2053));   // src/spi.v(275[8] 290[4])
    defparam i1700_4_lut.LUT_INIT = 16'hce0a;
    SB_LUT4 i1701_4_lut (.I0(tx_shift_reg[3]), .I1(tx_data_byte[4]), .I2(n3279), 
            .I3(n1728), .O(n2054));   // src/spi.v(275[8] 290[4])
    defparam i1701_4_lut.LUT_INIT = 16'hce0a;
    SB_LUT4 i1576_3_lut (.I0(tx_data_byte[0]), .I1(pc_data_rx[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n1929));   // src/top.v(748[8] 802[4])
    defparam i1576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1702_4_lut (.I0(tx_shift_reg[2]), .I1(tx_data_byte[3]), .I2(n3279), 
            .I3(n1728), .O(n2055));   // src/spi.v(275[8] 290[4])
    defparam i1702_4_lut.LUT_INIT = 16'hce0a;
    SB_LUT4 i1577_3_lut (.I0(\mem_LUT.mem_1_7 ), .I1(rx_buf_byte[7]), .I2(n4_adj_494), 
            .I3(GND_net), .O(n1930));   // src/fifo_quad_word_mod.v(448[73:76])
    defparam i1577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2889_4_lut (.I0(n1), .I1(fifo_read_cmd), .I2(wr_addr_r[1]), 
            .I3(rd_addr_r[1]), .O(n3275));
    defparam i2889_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i1703_3_lut (.I0(tx_data_byte[3]), .I1(pc_data_rx[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n2056));   // src/top.v(748[8] 802[4])
    defparam i1703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_581_788_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7), .I3(n2955), .O(n112)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_DFF reset_clk_counter_i3_582__i1 (.Q(reset_clk_counter[1]), .C(SLM_CLK_c), 
           .D(n2990));   // src/top.v(250[27:51])
    SB_LUT4 i1704_4_lut (.I0(tx_shift_reg[1]), .I1(tx_data_byte[2]), .I2(n3279), 
            .I3(n1728), .O(n2057));   // src/spi.v(275[8] 290[4])
    defparam i1704_4_lut.LUT_INIT = 16'hce0a;
    SB_IO DATA30_pad (.PACKAGE_PIN(DATA30), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA30_pad.PIN_TYPE = 6'b011001;
    defparam DATA30_pad.PULLUP = 1'b0;
    defparam DATA30_pad.NEG_TRIGGER = 1'b0;
    defparam DATA30_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA29_pad (.PACKAGE_PIN(DATA29), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA29_pad.PIN_TYPE = 6'b011001;
    defparam DATA29_pad.PULLUP = 1'b0;
    defparam DATA29_pad.NEG_TRIGGER = 1'b0;
    defparam DATA29_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA1_pad (.PACKAGE_PIN(DATA1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA1_pad.PIN_TYPE = 6'b011001;
    defparam DATA1_pad.PULLUP = 1'b0;
    defparam DATA1_pad.NEG_TRIGGER = 1'b0;
    defparam DATA1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA28_pad (.PACKAGE_PIN(DATA28), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA28_pad.PIN_TYPE = 6'b011001;
    defparam DATA28_pad.PULLUP = 1'b0;
    defparam DATA28_pad.NEG_TRIGGER = 1'b0;
    defparam DATA28_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA27_pad (.PACKAGE_PIN(DATA27), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA27_pad.PIN_TYPE = 6'b011001;
    defparam DATA27_pad.PULLUP = 1'b0;
    defparam DATA27_pad.NEG_TRIGGER = 1'b0;
    defparam DATA27_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA2_pad (.PACKAGE_PIN(DATA2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA2_pad.PIN_TYPE = 6'b011001;
    defparam DATA2_pad.PULLUP = 1'b0;
    defparam DATA2_pad.NEG_TRIGGER = 1'b0;
    defparam DATA2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA26_pad (.PACKAGE_PIN(DATA26), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA26_pad.PIN_TYPE = 6'b011001;
    defparam DATA26_pad.PULLUP = 1'b0;
    defparam DATA26_pad.NEG_TRIGGER = 1'b0;
    defparam DATA26_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA25_pad (.PACKAGE_PIN(DATA25), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA25_pad.PIN_TYPE = 6'b011001;
    defparam DATA25_pad.PULLUP = 1'b0;
    defparam DATA25_pad.NEG_TRIGGER = 1'b0;
    defparam DATA25_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA3_pad (.PACKAGE_PIN(DATA3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA3_pad.PIN_TYPE = 6'b011001;
    defparam DATA3_pad.PULLUP = 1'b0;
    defparam DATA3_pad.NEG_TRIGGER = 1'b0;
    defparam DATA3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA24_pad (.PACKAGE_PIN(DATA24), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA24_pad.PIN_TYPE = 6'b011001;
    defparam DATA24_pad.PULLUP = 1'b0;
    defparam DATA24_pad.NEG_TRIGGER = 1'b0;
    defparam DATA24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA23_pad (.PACKAGE_PIN(DATA23), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA23_pad.PIN_TYPE = 6'b011001;
    defparam DATA23_pad.PULLUP = 1'b0;
    defparam DATA23_pad.NEG_TRIGGER = 1'b0;
    defparam DATA23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA4_pad (.PACKAGE_PIN(DATA4), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA4_pad.PIN_TYPE = 6'b011001;
    defparam DATA4_pad.PULLUP = 1'b0;
    defparam DATA4_pad.NEG_TRIGGER = 1'b0;
    defparam DATA4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA22_pad (.PACKAGE_PIN(DATA22), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA22_pad.PIN_TYPE = 6'b011001;
    defparam DATA22_pad.PULLUP = 1'b0;
    defparam DATA22_pad.NEG_TRIGGER = 1'b0;
    defparam DATA22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA21_pad (.PACKAGE_PIN(DATA21), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA21_pad.PIN_TYPE = 6'b011001;
    defparam DATA21_pad.PULLUP = 1'b0;
    defparam DATA21_pad.NEG_TRIGGER = 1'b0;
    defparam DATA21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA5_pad (.PACKAGE_PIN(DATA5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA5_pad.PIN_TYPE = 6'b011001;
    defparam DATA5_pad.PULLUP = 1'b0;
    defparam DATA5_pad.NEG_TRIGGER = 1'b0;
    defparam DATA5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA20_pad (.PACKAGE_PIN(DATA20), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA20_pad.PIN_TYPE = 6'b011001;
    defparam DATA20_pad.PULLUP = 1'b0;
    defparam DATA20_pad.NEG_TRIGGER = 1'b0;
    defparam DATA20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA19_pad (.PACKAGE_PIN(DATA19), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA19_pad.PIN_TYPE = 6'b011001;
    defparam DATA19_pad.PULLUP = 1'b0;
    defparam DATA19_pad.NEG_TRIGGER = 1'b0;
    defparam DATA19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA6_pad (.PACKAGE_PIN(DATA6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA6_pad.PIN_TYPE = 6'b011001;
    defparam DATA6_pad.PULLUP = 1'b0;
    defparam DATA6_pad.NEG_TRIGGER = 1'b0;
    defparam DATA6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA18_pad (.PACKAGE_PIN(DATA18), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA18_pad.PIN_TYPE = 6'b011001;
    defparam DATA18_pad.PULLUP = 1'b0;
    defparam DATA18_pad.NEG_TRIGGER = 1'b0;
    defparam DATA18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA17_pad (.PACKAGE_PIN(DATA17), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA17_pad.PIN_TYPE = 6'b011001;
    defparam DATA17_pad.PULLUP = 1'b0;
    defparam DATA17_pad.NEG_TRIGGER = 1'b0;
    defparam DATA17_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA7_pad (.PACKAGE_PIN(DATA7), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA7_pad.PIN_TYPE = 6'b011001;
    defparam DATA7_pad.PULLUP = 1'b0;
    defparam DATA7_pad.NEG_TRIGGER = 1'b0;
    defparam DATA7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA16_pad (.PACKAGE_PIN(DATA16), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA16_pad.PIN_TYPE = 6'b011001;
    defparam DATA16_pad.PULLUP = 1'b0;
    defparam DATA16_pad.NEG_TRIGGER = 1'b0;
    defparam DATA16_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA15_pad (.PACKAGE_PIN(DATA15), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA15_pad.PIN_TYPE = 6'b011001;
    defparam DATA15_pad.PULLUP = 1'b0;
    defparam DATA15_pad.NEG_TRIGGER = 1'b0;
    defparam DATA15_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA8_pad (.PACKAGE_PIN(DATA8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA8_pad.PIN_TYPE = 6'b011001;
    defparam DATA8_pad.PULLUP = 1'b0;
    defparam DATA8_pad.NEG_TRIGGER = 1'b0;
    defparam DATA8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA14_pad (.PACKAGE_PIN(DATA14), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA14_pad.PIN_TYPE = 6'b011001;
    defparam DATA14_pad.PULLUP = 1'b0;
    defparam DATA14_pad.NEG_TRIGGER = 1'b0;
    defparam DATA14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA13_pad (.PACKAGE_PIN(DATA13), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA13_pad.PIN_TYPE = 6'b011001;
    defparam DATA13_pad.PULLUP = 1'b0;
    defparam DATA13_pad.NEG_TRIGGER = 1'b0;
    defparam DATA13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA12_pad (.PACKAGE_PIN(DATA12), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA12_pad.PIN_TYPE = 6'b011001;
    defparam DATA12_pad.PULLUP = 1'b0;
    defparam DATA12_pad.NEG_TRIGGER = 1'b0;
    defparam DATA12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA11_pad (.PACKAGE_PIN(DATA11), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA11_pad.PIN_TYPE = 6'b011001;
    defparam DATA11_pad.PULLUP = 1'b0;
    defparam DATA11_pad.NEG_TRIGGER = 1'b0;
    defparam DATA11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA9_pad (.PACKAGE_PIN(DATA9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA9_pad.PIN_TYPE = 6'b011001;
    defparam DATA9_pad.PULLUP = 1'b0;
    defparam DATA9_pad.NEG_TRIGGER = 1'b0;
    defparam DATA9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA10_pad (.PACKAGE_PIN(DATA10), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA10_pad.PIN_TYPE = 6'b011001;
    defparam DATA10_pad.PULLUP = 1'b0;
    defparam DATA10_pad.NEG_TRIGGER = 1'b0;
    defparam DATA10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_OE_pad (.PACKAGE_PIN(FT_OE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(FT_OE_c));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_OE_pad.PIN_TYPE = 6'b011001;
    defparam FT_OE_pad.PULLUP = 1'b0;
    defparam FT_OE_pad.NEG_TRIGGER = 1'b0;
    defparam FT_OE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_RD_pad (.PACKAGE_PIN(FT_RD), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(FT_RD_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_RD_pad.PIN_TYPE = 6'b011001;
    defparam FT_RD_pad.PULLUP = 1'b0;
    defparam FT_RD_pad.NEG_TRIGGER = 1'b0;
    defparam FT_RD_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_WR_pad (.PACKAGE_PIN(FT_WR), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_WR_pad.PIN_TYPE = 6'b101001;
    defparam FT_WR_pad.PULLUP = 1'b0;
    defparam FT_WR_pad.NEG_TRIGGER = 1'b0;
    defparam FT_WR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_SIWU_pad (.PACKAGE_PIN(FT_SIWU), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_SIWU_pad.PIN_TYPE = 6'b101001;
    defparam FT_SIWU_pad.PULLUP = 1'b0;
    defparam FT_SIWU_pad.NEG_TRIGGER = 1'b0;
    defparam FT_SIWU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_BE3_pad (.PACKAGE_PIN(FIFO_BE3), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_BE3_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_BE3_pad.PULLUP = 1'b0;
    defparam FIFO_BE3_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_BE3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_BE2_pad (.PACKAGE_PIN(FIFO_BE2), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_BE2_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_BE2_pad.PULLUP = 1'b0;
    defparam FIFO_BE2_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_BE2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1637_2_lut (.I0(spi_busy), .I1(spi_busy_prev), .I2(GND_net), 
            .I3(GND_net), .O(n1990));   // src/top.v(552[8] 558[4])
    defparam i1637_2_lut.LUT_INIT = 16'h4444;
    SB_IO FIFO_BE1_pad (.PACKAGE_PIN(FIFO_BE1), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_BE1_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_BE1_pad.PULLUP = 1'b0;
    defparam FIFO_BE1_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_BE1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_BE0_pad (.PACKAGE_PIN(FIFO_BE0), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_BE0_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_BE0_pad.PULLUP = 1'b0;
    defparam FIFO_BE0_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_BE0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1638_2_lut (.I0(is_tx_fifo_full_flag), .I1(spi_busy_falling_edge), 
            .I2(GND_net), .I3(GND_net), .O(n1991));   // src/top.v(560[8] 569[4])
    defparam i1638_2_lut.LUT_INIT = 16'h4444;
    SB_IO FIFO_D31_pad (.PACKAGE_PIN(FIFO_D31), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D31_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D31_pad.PULLUP = 1'b0;
    defparam FIFO_D31_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D31_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D30_pad (.PACKAGE_PIN(FIFO_D30), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D30_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D30_pad.PULLUP = 1'b0;
    defparam FIFO_D30_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D30_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1642_3_lut (.I0(tx_data_byte[7]), .I1(pc_data_rx[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n1995));   // src/top.v(748[8] 802[4])
    defparam i1642_3_lut.LUT_INIT = 16'hcaca;
    SB_IO FIFO_D29_pad (.PACKAGE_PIN(FIFO_D29), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D29_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D29_pad.PULLUP = 1'b0;
    defparam FIFO_D29_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D29_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY led_counter_581_788_add_4_9 (.CI(n2944), .I0(GND_net), .I1(n18), 
            .CO(n2945));
    SB_IO FIFO_D28_pad (.PACKAGE_PIN(FIFO_D28), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D28_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D28_pad.PULLUP = 1'b0;
    defparam FIFO_D28_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D28_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D27_pad (.PACKAGE_PIN(FIFO_D27), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D27_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D27_pad.PULLUP = 1'b0;
    defparam FIFO_D27_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D27_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D26_pad (.PACKAGE_PIN(FIFO_D26), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D26_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D26_pad.PULLUP = 1'b0;
    defparam FIFO_D26_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D26_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1641_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[7]), .I2(\mem_LUT.data_raw_r [7]), 
            .I3(n1795), .O(n1994));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i1641_4_lut.LUT_INIT = 16'h5044;
    SB_IO FIFO_D25_pad (.PACKAGE_PIN(FIFO_D25), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D25_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D25_pad.PULLUP = 1'b0;
    defparam FIFO_D25_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D25_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1643_3_lut (.I0(tx_data_byte[6]), .I1(pc_data_rx[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n1996));   // src/top.v(748[8] 802[4])
    defparam i1643_3_lut.LUT_INIT = 16'hcaca;
    SB_IO FIFO_D24_pad (.PACKAGE_PIN(FIFO_D24), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D24_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D24_pad.PULLUP = 1'b0;
    defparam FIFO_D24_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D23_pad (.PACKAGE_PIN(FIFO_D23), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D23_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D23_pad.PULLUP = 1'b0;
    defparam FIFO_D23_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1580_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[3]), .I2(\mem_LUT.data_raw_r [3]), 
            .I3(n1795), .O(n1933));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i1580_4_lut.LUT_INIT = 16'h5044;
    SB_IO FIFO_D22_pad (.PACKAGE_PIN(FIFO_D22), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D22_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D22_pad.PULLUP = 1'b0;
    defparam FIFO_D22_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1644_3_lut (.I0(tx_data_byte[5]), .I1(pc_data_rx[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n1997));   // src/top.v(748[8] 802[4])
    defparam i1644_3_lut.LUT_INIT = 16'hcaca;
    SB_IO FIFO_D21_pad (.PACKAGE_PIN(FIFO_D21), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D21_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D21_pad.PULLUP = 1'b0;
    defparam FIFO_D21_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D20_pad (.PACKAGE_PIN(FIFO_D20), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D20_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D20_pad.PULLUP = 1'b0;
    defparam FIFO_D20_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D19_pad (.PACKAGE_PIN(FIFO_D19), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D19_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D19_pad.PULLUP = 1'b0;
    defparam FIFO_D19_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 led_counter_581_788_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19), .I3(n2943), .O(n124)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_IO FIFO_D18_pad (.PACKAGE_PIN(FIFO_D18), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D18_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D18_pad.PULLUP = 1'b0;
    defparam FIFO_D18_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY led_counter_581_788_add_4_20 (.CI(n2955), .I0(GND_net), .I1(n7), 
            .CO(n2956));
    SB_IO FIFO_D17_pad (.PACKAGE_PIN(FIFO_D17), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D17_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D17_pad.PULLUP = 1'b0;
    defparam FIFO_D17_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D17_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1_2_lut_adj_19 (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_508));
    defparam i1_2_lut_adj_19.LUT_INIT = 16'h6666;
    SB_IO FIFO_D16_pad (.PACKAGE_PIN(FIFO_D16), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D16_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D16_pad.PULLUP = 1'b0;
    defparam FIFO_D16_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D16_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D15_pad (.PACKAGE_PIN(FIFO_D15), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D15_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D15_pad.PULLUP = 1'b0;
    defparam FIFO_D15_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D15_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D14_pad (.PACKAGE_PIN(FIFO_D14), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D14_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D14_pad.PULLUP = 1'b0;
    defparam FIFO_D14_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY led_counter_581_788_add_4_8 (.CI(n2943), .I0(GND_net), .I1(n19), 
            .CO(n2944));
    SB_IO FIFO_D13_pad (.PACKAGE_PIN(FIFO_D13), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D13_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D13_pad.PULLUP = 1'b0;
    defparam FIFO_D13_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D12_pad (.PACKAGE_PIN(FIFO_D12), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D12_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D12_pad.PULLUP = 1'b0;
    defparam FIFO_D12_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D11_pad (.PACKAGE_PIN(FIFO_D11), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D11_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D11_pad.PULLUP = 1'b0;
    defparam FIFO_D11_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D10_pad (.PACKAGE_PIN(FIFO_D10), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D10_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D10_pad.PULLUP = 1'b0;
    defparam FIFO_D10_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D9_pad (.PACKAGE_PIN(FIFO_D9), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D9_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D9_pad.PULLUP = 1'b0;
    defparam FIFO_D9_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1582_3_lut (.I0(\mem_LUT.mem_1_6 ), .I1(rx_buf_byte[6]), .I2(n4_adj_494), 
            .I3(GND_net), .O(n1935));   // src/fifo_quad_word_mod.v(448[73:76])
    defparam i1582_3_lut.LUT_INIT = 16'hcaca;
    SB_IO FIFO_D8_pad (.PACKAGE_PIN(FIFO_D8), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D8_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D8_pad.PULLUP = 1'b0;
    defparam FIFO_D8_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D7_pad (.PACKAGE_PIN(FIFO_D7), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D7_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D7_pad.PULLUP = 1'b0;
    defparam FIFO_D7_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D6_pad (.PACKAGE_PIN(FIFO_D6), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D6_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D6_pad.PULLUP = 1'b0;
    defparam FIFO_D6_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D5_pad (.PACKAGE_PIN(FIFO_D5), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D5_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D5_pad.PULLUP = 1'b0;
    defparam FIFO_D5_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D4_pad (.PACKAGE_PIN(FIFO_D4), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D4_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D4_pad.PULLUP = 1'b0;
    defparam FIFO_D4_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D3_pad (.PACKAGE_PIN(FIFO_D3), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D3_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D3_pad.PULLUP = 1'b0;
    defparam FIFO_D3_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D2_pad (.PACKAGE_PIN(FIFO_D2), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D2_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D2_pad.PULLUP = 1'b0;
    defparam FIFO_D2_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D1_pad (.PACKAGE_PIN(FIFO_D1), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D1_pad.PIN_TYPE = 6'b101001;
    defparam FIFO_D1_pad.PULLUP = 1'b0;
    defparam FIFO_D1_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_0_pad (.PACKAGE_PIN(DEBUG_0), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_0_c_24));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_0_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_0_pad.PULLUP = 1'b0;
    defparam DEBUG_0_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_1_pad (.PACKAGE_PIN(DEBUG_1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_1_c));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_1_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_1_pad.PULLUP = 1'b0;
    defparam DEBUG_1_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_2_pad (.PACKAGE_PIN(DEBUG_2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_2_c));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_2_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_2_pad.PULLUP = 1'b0;
    defparam DEBUG_2_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_3_pad (.PACKAGE_PIN(DEBUG_3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_3_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_3_pad.PULLUP = 1'b0;
    defparam DEBUG_3_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_5_pad (.PACKAGE_PIN(DEBUG_5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_5_c_c));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_5_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_5_pad.PULLUP = 1'b0;
    defparam DEBUG_5_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_6_pad (.PACKAGE_PIN(DEBUG_6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_6_c));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_6_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_6_pad.PULLUP = 1'b0;
    defparam DEBUG_6_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_8_pad (.PACKAGE_PIN(DEBUG_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_8_c_c));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_8_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_8_pad.PULLUP = 1'b0;
    defparam DEBUG_8_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_9_pad (.PACKAGE_PIN(DEBUG_9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_9_c_c));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_9_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_9_pad.PULLUP = 1'b0;
    defparam DEBUG_9_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CLK_pad (.PACKAGE_PIN(ICE_CLK), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CLK_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CLK_pad.PULLUP = 1'b0;
    defparam ICE_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CDONE_pad (.PACKAGE_PIN(ICE_CDONE), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CDONE_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CDONE_pad.PULLUP = 1'b0;
    defparam ICE_CDONE_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CDONE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CREST_pad (.PACKAGE_PIN(ICE_CREST), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CREST_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CREST_pad.PULLUP = 1'b0;
    defparam ICE_CREST_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CREST_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_SYSCLK_pad (.PACKAGE_PIN(ICE_SYSCLK), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ICE_SYSCLK_c));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_SYSCLK_pad.PIN_TYPE = 6'b000001;
    defparam ICE_SYSCLK_pad.PULLUP = 1'b0;
    defparam ICE_SYSCLK_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_SYSCLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UART_RX_pad (.PACKAGE_PIN(UART_RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(UART_RX_c)) /* synthesis IO_FF_IN=TRUE */ ;   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UART_RX_pad.PIN_TYPE = 6'b000001;
    defparam UART_RX_pad.PULLUP = 1'b0;
    defparam UART_RX_pad.NEG_TRIGGER = 1'b0;
    defparam UART_RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_5_c_pad (.PACKAGE_PIN(SOUT), .OUTPUT_ENABLE(VCC_net), .D_IN_0(DEBUG_5_c_c));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_5_c_pad.PIN_TYPE = 6'b000001;
    defparam DEBUG_5_c_pad.PULLUP = 1'b0;
    defparam DEBUG_5_c_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_5_c_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_9_c_pad (.PACKAGE_PIN(FR_RXF), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(DEBUG_9_c_c));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_9_c_pad.PIN_TYPE = 6'b000001;
    defparam DEBUG_9_c_pad.PULLUP = 1'b0;
    defparam DEBUG_9_c_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_9_c_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO FIFO_CLK_pad (.PACKAGE_PIN(FIFO_CLK), .OUTPUT_ENABLE(VCC_net), 
            .GLOBAL_BUFFER_OUTPUT(FIFO_CLK_c));   // src/top.v(84[12:20])
    defparam FIFO_CLK_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_CLK_pad.PULLUP = 1'b0;
    defparam FIFO_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_8_c_pad (.PACKAGE_PIN(FIFO_D0), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(DEBUG_8_c_c));   // C:/lscc/iCEcube2/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_8_c_pad.PIN_TYPE = 6'b000001;
    defparam DEBUG_8_c_pad.PULLUP = 1'b0;
    defparam DEBUG_8_c_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_8_c_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 led_counter_581_788_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20), .I3(n2942), .O(n125)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_581_788_add_4_7 (.CI(n2942), .I0(GND_net), .I1(n20), 
            .CO(n2943));
    SB_LUT4 led_counter_581_788_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_501), .I3(n2954), .O(n113)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 led_counter_581_788_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21), .I3(n2941), .O(n126)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_581_788_add_4_19 (.CI(n2954), .I0(GND_net), .I1(n8_adj_501), 
            .CO(n2955));
    SB_CARRY led_counter_581_788_add_4_6 (.CI(n2941), .I0(GND_net), .I1(n21), 
            .CO(n2942));
    SB_LUT4 led_counter_581_788_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9), .I3(n2953), .O(n114)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut (.I0(reset_all_w), .I1(n15_adj_509), .I2(wr_fifo_en_w), 
            .I3(n2968), .O(n3118));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut.LUT_INIT = 16'h5444;
    SB_LUT4 led_counter_581_788_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22), .I3(n2940), .O(n127)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_581_788_add_4_18 (.CI(n2953), .I0(GND_net), .I1(n9), 
            .CO(n2954));
    SB_CARRY led_counter_581_788_add_4_5 (.CI(n2940), .I0(GND_net), .I1(n22), 
            .CO(n2941));
    SB_DFF start_tx_206 (.Q(r_SM_Main_2__N_187[0]), .C(SLM_CLK_c), .D(n2010));   // src/top.v(581[8] 599[4])
    SB_LUT4 led_counter_581_788_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23), .I3(n2939), .O(n128)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1586_3_lut (.I0(\mem_LUT.mem_1_5 ), .I1(rx_buf_byte[5]), .I2(n4_adj_494), 
            .I3(GND_net), .O(n1939));   // src/fifo_quad_word_mod.v(448[73:76])
    defparam i1586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1705_3_lut (.I0(tx_data_byte[2]), .I1(pc_data_rx[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n2058));   // src/top.v(748[8] 802[4])
    defparam i1705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_581_788_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10), .I3(n2952), .O(n115)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1645_3_lut (.I0(tx_data_byte[4]), .I1(pc_data_rx[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n1998));   // src/top.v(748[8] 802[4])
    defparam i1645_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_581_788_add_4_4 (.CI(n2939), .I0(GND_net), .I1(n23), 
            .CO(n2940));
    SB_CARRY led_counter_581_788_add_4_17 (.CI(n2952), .I0(GND_net), .I1(n10), 
            .CO(n2953));
    SB_LUT4 led_counter_581_788_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11), .I3(n2951), .O(n116)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 led_counter_581_788_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24), .I3(n2938), .O(n129)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_581_788_add_4_3 (.CI(n2938), .I0(GND_net), .I1(n24), 
            .CO(n2939));
    SB_LUT4 i1706_4_lut (.I0(tx_shift_reg[0]), .I1(tx_data_byte[1]), .I2(n3279), 
            .I3(n1728), .O(n2059));   // src/spi.v(275[8] 290[4])
    defparam i1706_4_lut.LUT_INIT = 16'hce0a;
    SB_CARRY led_counter_581_788_add_4_16 (.CI(n2951), .I0(GND_net), .I1(n11), 
            .CO(n2952));
    SB_LUT4 led_counter_581_788_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12), .I3(n2950), .O(n117)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1646_3_lut (.I0(tx_addr_byte[7]), .I1(tx_data_byte[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n1999));   // src/top.v(748[8] 802[4])
    defparam i1646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_581_788_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25), .I3(VCC_net), .O(n130)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_108[2]), 
            .I3(r_SM_Main[0]), .O(n1764));   // src/uart_rx.v(49[10] 144[8])
    defparam i13_3_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i1707_3_lut (.I0(r_Tx_Data[7]), .I1(fifo_temp_output[7]), .I2(n1636), 
            .I3(GND_net), .O(n2060));   // src/uart_tx.v(38[10] 141[8])
    defparam i1707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_108[2]), 
            .I3(r_SM_Main[0]), .O(n3250));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_DFF reset_clk_counter_i3_582__i2 (.Q(reset_clk_counter[2]), .C(SLM_CLK_c), 
           .D(n2992));   // src/top.v(250[27:51])
    SB_DFF reset_clk_counter_i3_582__i3 (.Q(reset_clk_counter[3]), .C(SLM_CLK_c), 
           .D(n2994));   // src/top.v(250[27:51])
    SB_DFF tx_addr_byte_r_i0_i1 (.Q(tx_addr_byte[1]), .C(SLM_CLK_c), .D(n2005));   // src/top.v(748[8] 802[4])
    SB_DFF tx_addr_byte_r_i0_i2 (.Q(tx_addr_byte[2]), .C(SLM_CLK_c), .D(n2004));   // src/top.v(748[8] 802[4])
    SB_DFF tx_addr_byte_r_i0_i3 (.Q(tx_addr_byte[3]), .C(SLM_CLK_c), .D(n2003));   // src/top.v(748[8] 802[4])
    SB_DFF tx_addr_byte_r_i0_i4 (.Q(tx_addr_byte[4]), .C(SLM_CLK_c), .D(n2002));   // src/top.v(748[8] 802[4])
    SB_DFF tx_addr_byte_r_i0_i5 (.Q(tx_addr_byte[5]), .C(SLM_CLK_c), .D(n2001));   // src/top.v(748[8] 802[4])
    SB_DFF tx_addr_byte_r_i0_i6 (.Q(tx_addr_byte[6]), .C(SLM_CLK_c), .D(n2000));   // src/top.v(748[8] 802[4])
    SB_DFF tx_addr_byte_r_i0_i7 (.Q(tx_addr_byte[7]), .C(SLM_CLK_c), .D(n1999));   // src/top.v(748[8] 802[4])
    SB_DFF tx_data_byte_r_i0_i4 (.Q(tx_data_byte[4]), .C(SLM_CLK_c), .D(n1998));   // src/top.v(748[8] 802[4])
    SB_DFF tx_data_byte_r_i0_i5 (.Q(tx_data_byte[5]), .C(SLM_CLK_c), .D(n1997));   // src/top.v(748[8] 802[4])
    SB_DFF tx_data_byte_r_i0_i6 (.Q(tx_data_byte[6]), .C(SLM_CLK_c), .D(n1996));   // src/top.v(748[8] 802[4])
    SB_DFF tx_data_byte_r_i0_i7 (.Q(tx_data_byte[7]), .C(SLM_CLK_c), .D(n1995));   // src/top.v(748[8] 802[4])
    SB_DFF fifo_write_cmd_204 (.Q(fifo_write_cmd), .C(SLM_CLK_c), .D(n1991));   // src/top.v(560[8] 569[4])
    SB_DFF spi_busy_falling_edge_202 (.Q(spi_busy_falling_edge), .C(SLM_CLK_c), 
           .D(n1990));   // src/top.v(552[8] 558[4])
    SB_LUT4 i1647_3_lut (.I0(tx_addr_byte[6]), .I1(tx_data_byte[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n2000));   // src/top.v(748[8] 802[4])
    defparam i1647_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_data_byte_r_i0_i0 (.Q(tx_data_byte[0]), .C(SLM_CLK_c), .D(n1929));   // src/top.v(748[8] 802[4])
    SB_DFF uart_rx_complete_rising_edge_207 (.Q(uart_rx_complete_rising_edge), 
           .C(SLM_CLK_c), .D(n1988));   // src/top.v(739[8] 745[4])
    SB_CARRY led_counter_581_788_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(n25), 
            .CO(n2938));
    SB_LUT4 i1648_3_lut (.I0(tx_addr_byte[5]), .I1(tx_data_byte[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n2001));   // src/top.v(748[8] 802[4])
    defparam i1648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1649_3_lut (.I0(tx_addr_byte[4]), .I1(tx_data_byte[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n2002));   // src/top.v(748[8] 802[4])
    defparam i1649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1650_3_lut (.I0(tx_addr_byte[3]), .I1(tx_data_byte[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n2003));   // src/top.v(748[8] 802[4])
    defparam i1650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1608_3_lut (.I0(tx_addr_byte[0]), .I1(tx_data_byte[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n1961));   // src/top.v(748[8] 802[4])
    defparam i1608_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_581_788_add_4_15 (.CI(n2950), .I0(GND_net), .I1(n12), 
            .CO(n2951));
    SB_LUT4 i1651_3_lut (.I0(tx_addr_byte[2]), .I1(tx_data_byte[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n2004));   // src/top.v(748[8] 802[4])
    defparam i1651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1652_3_lut (.I0(tx_addr_byte[1]), .I1(tx_data_byte[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n2005));   // src/top.v(748[8] 802[4])
    defparam i1652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_20 (.I0(DEBUG_5_c_c), .I1(n3279), .I2(GND_net), 
            .I3(GND_net), .O(n3178));   // src/spi.v(299[8] 313[4])
    defparam i1_2_lut_adj_20.LUT_INIT = 16'h2222;
    SB_LUT4 led_counter_581_788_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13), .I3(n2949), .O(n118)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_DFF debug_check_211 (.Q(DEBUG_2_c), .C(SLM_CLK_c), .D(n1982));   // src/top.v(748[8] 802[4])
    SB_CARRY led_counter_581_788_add_4_14 (.CI(n2949), .I0(GND_net), .I1(n13), 
            .CO(n2950));
    GND i1 (.Y(GND_net));
    SB_DFF FT_OE_r_200 (.Q(FT_OE_c), .C(FIFO_CLK_c), .D(DEBUG_9_c_c));   // src/top.v(289[8] 303[6])
    SB_LUT4 i1708_3_lut (.I0(r_Tx_Data[6]), .I1(fifo_temp_output[6]), .I2(n1636), 
            .I3(GND_net), .O(n2061));   // src/uart_tx.v(38[10] 141[8])
    defparam i1708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1709_3_lut (.I0(r_Tx_Data[5]), .I1(fifo_temp_output[5]), .I2(n1636), 
            .I3(GND_net), .O(n2062));   // src/uart_tx.v(38[10] 141[8])
    defparam i1709_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_581_788_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14), .I3(n2948), .O(n119)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_581_788_add_4_13 (.CI(n2948), .I0(GND_net), .I1(n14), 
            .CO(n2949));
    SB_LUT4 led_counter_581_788_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15), .I3(n2947), .O(n120)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_581_788_add_4_12 (.CI(n2947), .I0(GND_net), .I1(n15), 
            .CO(n2948));
    SB_LUT4 led_counter_581_788_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16), .I3(n2946), .O(n121)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 led_counter_581_788_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(DEBUG_0_c_24), .I3(n2961), .O(n106)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 led_counter_581_788_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n2_adj_503), .I3(n2960), .O(n107)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_581_788_add_4_25 (.CI(n2960), .I0(GND_net), .I1(n2_adj_503), 
            .CO(n2961));
    SB_LUT4 led_counter_581_788_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3), .I3(n2959), .O(n108)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_581_788_add_4_24 (.CI(n2959), .I0(GND_net), .I1(n3), 
            .CO(n2960));
    SB_LUT4 led_counter_581_788_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_502), .I3(n2958), .O(n109)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_581_788_add_4_23 (.CI(n2958), .I0(GND_net), .I1(n4_adj_502), 
            .CO(n2959));
    SB_LUT4 led_counter_581_788_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5), .I3(n2957), .O(n110)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_581_788_add_4_22 (.CI(n2957), .I0(GND_net), .I1(n5), 
            .CO(n2958));
    SB_LUT4 led_counter_581_788_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6), .I3(n2956), .O(n111)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_581_788_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1591_3_lut (.I0(\mem_LUT.mem_1_4 ), .I1(rx_buf_byte[4]), .I2(n4_adj_494), 
            .I3(GND_net), .O(n1944));   // src/fifo_quad_word_mod.v(448[73:76])
    defparam i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1592_3_lut (.I0(\mem_LUT.mem_1_3 ), .I1(rx_buf_byte[3]), .I2(n4_adj_494), 
            .I3(GND_net), .O(n1945));   // src/fifo_quad_word_mod.v(448[73:76])
    defparam i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1609_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[1]), .I2(n4_adj_500), 
            .I3(n1754), .O(n1962));   // src/uart_rx.v(49[10] 144[8])
    defparam i1609_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1597_3_lut (.I0(r_Tx_Data[0]), .I1(fifo_temp_output[0]), .I2(n1636), 
            .I3(GND_net), .O(n1950));   // src/uart_tx.v(38[10] 141[8])
    defparam i1597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1598_3_lut (.I0(\mem_LUT.mem_1_2 ), .I1(rx_buf_byte[2]), .I2(n4_adj_494), 
            .I3(GND_net), .O(n1951));   // src/fifo_quad_word_mod.v(448[73:76])
    defparam i1598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1601_3_lut (.I0(\mem_LUT.mem_1_1 ), .I1(rx_buf_byte[1]), .I2(n4_adj_494), 
            .I3(GND_net), .O(n1954));   // src/fifo_quad_word_mod.v(448[73:76])
    defparam i1601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1711_3_lut (.I0(r_Tx_Data[4]), .I1(fifo_temp_output[4]), .I2(n1636), 
            .I3(GND_net), .O(n2064));   // src/uart_tx.v(38[10] 141[8])
    defparam i1711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1712_3_lut (.I0(r_Tx_Data[3]), .I1(fifo_temp_output[3]), .I2(n1636), 
            .I3(GND_net), .O(n2065));   // src/uart_tx.v(38[10] 141[8])
    defparam i1712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1610_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[2]), .I2(n4_adj_504), 
            .I3(n1750), .O(n1963));   // src/uart_rx.v(49[10] 144[8])
    defparam i1610_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1603_3_lut (.I0(rx_buf_byte[0]), .I1(rx_shift_reg[1]), .I2(rx_shift_reg_15__N_319), 
            .I3(GND_net), .O(n1956));   // src/spi.v(299[8] 313[4])
    defparam i1603_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1713_3_lut (.I0(r_Tx_Data[2]), .I1(fifo_temp_output[2]), .I2(n1636), 
            .I3(GND_net), .O(n2066));   // src/uart_tx.v(38[10] 141[8])
    defparam i1713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1604_3_lut (.I0(\mem_LUT.mem_1_0 ), .I1(rx_buf_byte[0]), .I2(n4_adj_494), 
            .I3(GND_net), .O(n1957));   // src/fifo_quad_word_mod.v(448[73:76])
    defparam i1604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2550_2_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_505));   // src/top.v(250[27:51])
    defparam i2550_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1714_3_lut (.I0(r_Tx_Data[1]), .I1(fifo_temp_output[1]), .I2(n1636), 
            .I3(GND_net), .O(n2067));   // src/uart_tx.v(38[10] 141[8])
    defparam i1714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1715_3_lut (.I0(tx_data_byte[1]), .I1(pc_data_rx[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n2068));   // src/top.v(748[8] 802[4])
    defparam i1715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_21 (.I0(rx_shift_reg[0]), .I1(n3279), .I2(GND_net), 
            .I3(GND_net), .O(n3180));   // src/spi.v(299[8] 313[4])
    defparam i1_2_lut_adj_21.LUT_INIT = 16'h2222;
    SB_LUT4 i1672_3_lut (.I0(rx_buf_byte[7]), .I1(rx_shift_reg[8]), .I2(rx_shift_reg_15__N_319), 
            .I3(GND_net), .O(n2025));   // src/spi.v(299[8] 313[4])
    defparam i1672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1663_4_lut (.I0(n3293), .I1(r_Bit_Index[0]), .I2(n2540), 
            .I3(r_SM_Main[1]), .O(n2016));   // src/uart_rx.v(49[10] 144[8])
    defparam i1663_4_lut.LUT_INIT = 16'h4644;
    SB_LUT4 i1676_3_lut (.I0(rx_buf_byte[6]), .I1(rx_shift_reg[7]), .I2(rx_shift_reg_15__N_319), 
            .I3(GND_net), .O(n2029));   // src/spi.v(299[8] 313[4])
    defparam i1676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_22 (.I0(start_transfer_edge), .I1(start_transfer_prev), 
            .I2(n5_adj_507), .I3(DEBUG_2_c), .O(n3148));   // src/spi.v(73[8] 82[4])
    defparam i1_4_lut_adj_22.LUT_INIT = 16'hb3a0;
    SB_LUT4 i1677_3_lut (.I0(rx_buf_byte[5]), .I1(rx_shift_reg[6]), .I2(rx_shift_reg_15__N_319), 
            .I3(GND_net), .O(n2030));   // src/spi.v(299[8] 313[4])
    defparam i1677_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1678_3_lut (.I0(rx_buf_byte[4]), .I1(rx_shift_reg[5]), .I2(rx_shift_reg_15__N_319), 
            .I3(GND_net), .O(n2031));   // src/spi.v(299[8] 313[4])
    defparam i1678_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1028_2_lut_3_lut_4_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(reset_all_w), .I3(wr_addr_r[0]), .O(n8));
    defparam i1028_2_lut_3_lut_4_lut.LUT_INIT = 16'h0df2;
    SB_LUT4 i1_3_lut_4_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(wr_addr_r[0]), .I3(rd_addr_r[0]), .O(n4_adj_511));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0220;
    SB_LUT4 i1679_3_lut (.I0(rx_buf_byte[3]), .I1(rx_shift_reg[4]), .I2(rx_shift_reg_15__N_319), 
            .I3(GND_net), .O(n2032));   // src/spi.v(299[8] 313[4])
    defparam i1679_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1680_3_lut (.I0(rx_buf_byte[2]), .I1(rx_shift_reg[3]), .I2(rx_shift_reg_15__N_319), 
            .I3(GND_net), .O(n2033));   // src/spi.v(299[8] 313[4])
    defparam i1680_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1681_3_lut (.I0(rx_buf_byte[1]), .I1(rx_shift_reg[2]), .I2(rx_shift_reg_15__N_319), 
            .I3(GND_net), .O(n2034));   // src/spi.v(299[8] 313[4])
    defparam i1681_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1682_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[0]), .I2(n4_adj_500), 
            .I3(n1750), .O(n2035));   // src/uart_rx.v(49[10] 144[8])
    defparam i1682_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1660_3_lut (.I0(n1898), .I1(r_Bit_Index_adj_514[0]), .I2(n1819), 
            .I3(GND_net), .O(n2013));   // src/uart_tx.v(38[10] 141[8])
    defparam i1660_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i1_2_lut_adj_23 (.I0(rx_shift_reg[1]), .I1(n3279), .I2(GND_net), 
            .I3(GND_net), .O(n3184));   // src/spi.v(299[8] 313[4])
    defparam i1_2_lut_adj_23.LUT_INIT = 16'h2222;
    SB_LUT4 i1683_4_lut (.I0(tx_shift_reg[13]), .I1(tx_addr_byte[6]), .I2(n3279), 
            .I3(n1728), .O(n2036));   // src/spi.v(275[8] 290[4])
    defparam i1683_4_lut.LUT_INIT = 16'hce0a;
    SB_LUT4 i1684_4_lut (.I0(tx_shift_reg[12]), .I1(tx_addr_byte[5]), .I2(n3279), 
            .I3(n1728), .O(n2037));   // src/spi.v(275[8] 290[4])
    defparam i1684_4_lut.LUT_INIT = 16'hce0a;
    SB_LUT4 i1685_4_lut (.I0(tx_shift_reg[11]), .I1(tx_addr_byte[4]), .I2(n3279), 
            .I3(n1728), .O(n2038));   // src/spi.v(275[8] 290[4])
    defparam i1685_4_lut.LUT_INIT = 16'hce0a;
    SB_LUT4 i1686_4_lut (.I0(tx_shift_reg[10]), .I1(tx_addr_byte[3]), .I2(n3279), 
            .I3(n1728), .O(n2039));   // src/spi.v(275[8] 290[4])
    defparam i1686_4_lut.LUT_INIT = 16'hce0a;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(reset_clk_counter[1]), .I1(reset_all_w_N_61), 
            .I2(reset_clk_counter[0]), .I3(reset_clk_counter[2]), .O(n2992));   // src/top.v(250[27:51])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfb04;
    SB_LUT4 i1_4_lut_4_lut (.I0(is_tx_fifo_full_flag), .I1(n3275), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_509));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1687_4_lut (.I0(tx_shift_reg[9]), .I1(tx_addr_byte[2]), .I2(n3279), 
            .I3(n1728), .O(n2040));   // src/spi.v(275[8] 290[4])
    defparam i1687_4_lut.LUT_INIT = 16'hce0a;
    SB_LUT4 i1688_4_lut (.I0(tx_shift_reg[8]), .I1(tx_addr_byte[1]), .I2(n3279), 
            .I3(n1728), .O(n2041));   // src/spi.v(275[8] 290[4])
    defparam i1688_4_lut.LUT_INIT = 16'hce0a;
    SB_LUT4 i1689_4_lut (.I0(tx_shift_reg[7]), .I1(tx_addr_byte[0]), .I2(n3279), 
            .I3(n1728), .O(n2042));   // src/spi.v(275[8] 290[4])
    defparam i1689_4_lut.LUT_INIT = 16'hce0a;
    SB_LUT4 i1016_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n1285));   // src/top.v(748[8] 802[4])
    defparam i1016_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_24 (.I0(rx_shift_reg[2]), .I1(n3279), .I2(GND_net), 
            .I3(GND_net), .O(n3188));   // src/spi.v(299[8] 313[4])
    defparam i1_2_lut_adj_24.LUT_INIT = 16'h2222;
    SB_LUT4 i1690_4_lut (.I0(tx_shift_reg[6]), .I1(tx_data_byte[7]), .I2(n3279), 
            .I3(n1728), .O(n2043));   // src/spi.v(275[8] 290[4])
    defparam i1690_4_lut.LUT_INIT = 16'hce0a;
    SB_LUT4 i1691_3_lut (.I0(\mem_LUT.mem_3_0 ), .I1(rx_buf_byte[0]), .I2(n2), 
            .I3(GND_net), .O(n2044));   // src/fifo_quad_word_mod.v(448[73:76])
    defparam i1691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1692_3_lut (.I0(\mem_LUT.mem_3_1 ), .I1(rx_buf_byte[1]), .I2(n2), 
            .I3(GND_net), .O(n2045));   // src/fifo_quad_word_mod.v(448[73:76])
    defparam i1692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1693_3_lut (.I0(\mem_LUT.mem_3_2 ), .I1(rx_buf_byte[2]), .I2(n2), 
            .I3(GND_net), .O(n2046));   // src/fifo_quad_word_mod.v(448[73:76])
    defparam i1693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1694_3_lut (.I0(\mem_LUT.mem_3_3 ), .I1(rx_buf_byte[3]), .I2(n2), 
            .I3(GND_net), .O(n2047));   // src/fifo_quad_word_mod.v(448[73:76])
    defparam i1694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_25 (.I0(rx_shift_reg[3]), .I1(n3279), .I2(GND_net), 
            .I3(GND_net), .O(n3190));   // src/spi.v(299[8] 313[4])
    defparam i1_2_lut_adj_25.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_26 (.I0(rx_shift_reg[7]), .I1(n3279), .I2(GND_net), 
            .I3(GND_net), .O(n3212));   // src/spi.v(299[8] 313[4])
    defparam i1_2_lut_adj_26.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_27 (.I0(rx_shift_reg[4]), .I1(n3279), .I2(GND_net), 
            .I3(GND_net), .O(n3198));   // src/spi.v(299[8] 313[4])
    defparam i1_2_lut_adj_27.LUT_INIT = 16'h2222;
    SB_LUT4 i1656_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[0]), 
            .I2(\mem_LUT.data_raw_r [0]), .I3(n1795), .O(n2009));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i1656_4_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i2974_2_lut (.I0(is_fifo_empty_flag), .I1(tx_uart_active_flag), 
            .I2(GND_net), .I3(GND_net), .O(start_tx_N_71));
    defparam i2974_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_512[2]), .I1(r_SM_Main_2__N_184[1]), 
            .I2(r_SM_Main_adj_512[0]), .I3(r_SM_Main_adj_512[1]), .O(n3439));   // src/uart_tx.v(38[10] 141[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i1723_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[2]), 
            .I2(\mem_LUT.data_raw_r [2]), .I3(n1795), .O(n2076));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i1723_4_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i1720_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[1]), 
            .I2(\mem_LUT.data_raw_r [1]), .I3(n1795), .O(n2073));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i1720_4_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i1589_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[4]), .I2(\mem_LUT.data_raw_r [4]), 
            .I3(n1795), .O(n1942));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i1589_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i1_2_lut_3_lut (.I0(reset_clk_counter[1]), .I1(reset_all_w_N_61), 
            .I2(reset_clk_counter[0]), .I3(GND_net), .O(n2990));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'ha6a6;
    SB_LUT4 i1657_3_lut_4_lut (.I0(r_SM_Main_2__N_187[0]), .I1(fifo_read_cmd), 
            .I2(is_fifo_empty_flag), .I3(tx_uart_active_flag), .O(n2010));   // src/top.v(581[8] 599[4])
    defparam i1657_3_lut_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1596_4_lut_4_lut (.I0(tx_uart_active_flag), .I1(r_SM_Main_adj_512[1]), 
            .I2(r_SM_Main_adj_512[2]), .I3(n4), .O(n1949));   // src/uart_tx.v(38[10] 141[8])
    defparam i1596_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i1618_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[6]), .I2(\mem_LUT.data_raw_r [6]), 
            .I3(n1795), .O(n1971));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i1618_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_28 (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(reset_all_w), .I3(rd_fifo_en_prev_r), .O(n1795));
    defparam i1_2_lut_3_lut_4_lut_adj_28.LUT_INIT = 16'hfff2;
    SB_LUT4 i1630_2_lut_3_lut (.I0(reset_all_w), .I1(fifo_read_cmd), .I2(is_fifo_empty_flag), 
            .I3(GND_net), .O(n1983));   // src/fifo_quad_word_mod.v(353[29] 363[32])
    defparam i1630_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i529_4_lut (.I0(state_reg[1]), .I1(state_next_2__N_312), .I2(state_reg[2]), 
            .I3(state_reg[0]), .O(n883));   // src/spi.v(132[10:19])
    defparam i529_4_lut.LUT_INIT = 16'h4a40;
    SB_LUT4 i1027_2_lut_3_lut_4_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(reset_all_w), .I3(rd_addr_r[0]), .O(n8_adj_499));
    defparam i1027_2_lut_3_lut_4_lut.LUT_INIT = 16'h0df2;
    SB_LUT4 i1_3_lut_4_lut_adj_29 (.I0(reset_clk_counter[1]), .I1(n2_adj_505), 
            .I2(reset_clk_counter[2]), .I3(reset_clk_counter[3]), .O(n2994));   // src/top.v(250[27:51])
    defparam i1_3_lut_4_lut_adj_29.LUT_INIT = 16'hfe01;
    SB_LUT4 i1_4_lut_adj_30 (.I0(reset_all_w), .I1(n3289), .I2(n24_adj_510), 
            .I3(n4_adj_511), .O(n3239));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_adj_30.LUT_INIT = 16'hfbfa;
    SB_LUT4 i1595_4_lut_4_lut (.I0(wr_fifo_en_w), .I1(reset_all_w), .I2(wr_addr_p1_w[2]), 
            .I3(wr_addr_r[2]), .O(n1948));
    defparam i1595_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i1615_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[5]), .I2(\mem_LUT.data_raw_r [5]), 
            .I3(n1795), .O(n1968));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i1615_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i1_4_lut_adj_31 (.I0(rd_addr_r[1]), .I1(rd_addr_r[0]), .I2(wr_addr_r[1]), 
            .I3(wr_addr_r[0]), .O(n32));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_adj_31.LUT_INIT = 16'h8421;
    SB_LUT4 i1_3_lut (.I0(is_fifo_empty_flag), .I1(fifo_write_cmd), .I2(n32), 
            .I3(GND_net), .O(n24_adj_510));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i2902_4_lut (.I0(rd_addr_p1_w[2]), .I1(n3448), .I2(wr_addr_r[2]), 
            .I3(wr_addr_r[1]), .O(n3289));
    defparam i2902_4_lut.LUT_INIT = 16'h7bde;
    \uart_rx(CLKS_PER_BIT=434)  pc_rx (.r_Rx_Data(r_Rx_Data), .SLM_CLK_c(SLM_CLK_c), 
            .n1965(n1965), .pc_data_rx({pc_data_rx}), .\r_SM_Main_2__N_108[2] (r_SM_Main_2__N_108[2]), 
            .GND_net(GND_net), .n3250(n3250), .r_SM_Main({r_SM_Main}), 
            .n2016(n2016), .r_Bit_Index({Open_0, Open_1, r_Bit_Index[0]}), 
            .n1963(n1963), .n1962(n1962), .DEBUG_1_c(DEBUG_1_c), .n4(n4_adj_506), 
            .n3293(n3293), .n1747(n1747), .n2035(n2035), .uart_rx_complete_prev(uart_rx_complete_prev), 
            .n1988(n1988), .n2540(n2540), .VCC_net(VCC_net), .n1975(n1975), 
            .n1974(n1974), .n1973(n1973), .n1972(n1972), .UART_RX_c(UART_RX_c), 
            .n1764(n1764), .n4_adj_3(n4_adj_500), .n1750(n1750), .n1754(n1754), 
            .n4_adj_4(n4_adj_504)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(381[42] 386[3])
    SB_LUT4 i1585_4_lut_4_lut_4_lut (.I0(wr_fifo_en_w), .I1(reset_all_w), 
            .I2(wr_addr_r[0]), .I3(wr_addr_r[1]), .O(n1938));
    defparam i1585_4_lut_4_lut_4_lut.LUT_INIT = 16'h1320;
    clock clock_inst (.GND_net(GND_net), .VCC_net(VCC_net), .ICE_SYSCLK_c(ICE_SYSCLK_c), 
          .pll_clk_unbuf(pll_clk_unbuf)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(214[7] 219[3])
    SB_LUT4 i3_4_lut (.I0(reset_clk_counter[0]), .I1(reset_clk_counter[2]), 
            .I2(reset_clk_counter[3]), .I3(reset_clk_counter[1]), .O(reset_all_w_N_61));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    FIFO_Quad_Word tx_fifo (.rd_fifo_en_w(rd_fifo_en_w), .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r [0]), 
            .SLM_CLK_c(SLM_CLK_c), .n3239(n3239), .is_fifo_empty_flag(is_fifo_empty_flag), 
            .n1968(n1968), .\fifo_temp_output[5] (fifo_temp_output[5]), 
            .rd_addr_r({rd_addr_r}), .\mem_LUT.mem_3_5 (\mem_LUT.mem_3_5 ), 
            .n1971(n1971), .\fifo_temp_output[6] (fifo_temp_output[6]), 
            .\mem_LUT.mem_1_5 (\mem_LUT.mem_1_5 ), .n1978(n1978), .n1981(n1981), 
            .n3118(n3118), .is_tx_fifo_full_flag(is_tx_fifo_full_flag), 
            .n1933(n1933), .\fifo_temp_output[3] (fifo_temp_output[3]), 
            .n1994(n1994), .\fifo_temp_output[7] (fifo_temp_output[7]), 
            .n1938(n1938), .wr_addr_r({wr_addr_r}), .n1942(n1942), .\fifo_temp_output[4] (fifo_temp_output[4]), 
            .n8(n8), .reset_all_w(reset_all_w), .n1948(n1948), .n8_adj_2(n8_adj_499), 
            .n2009(n2009), .\fifo_temp_output[0] (fifo_temp_output[0]), 
            .fifo_write_cmd(fifo_write_cmd), .wr_fifo_en_w(wr_fifo_en_w), 
            .GND_net(GND_net), .n2076(n2076), .VCC_net(VCC_net), .\fifo_temp_output[2] (fifo_temp_output[2]), 
            .n2073(n2073), .\fifo_temp_output[1] (fifo_temp_output[1]), 
            .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r [7]), .n1(n1), 
            .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r [6]), .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r [5]), 
            .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r [4]), .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r [3]), 
            .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r [2]), .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r [1]), 
            .n2051(n2051), .\mem_LUT.mem_3_7 (\mem_LUT.mem_3_7 ), .n2050(n2050), 
            .\mem_LUT.mem_3_6 (\mem_LUT.mem_3_6 ), .\mem_LUT.mem_3_4 (\mem_LUT.mem_3_4 ), 
            .\mem_LUT.mem_1_4 (\mem_LUT.mem_1_4 ), .n2049(n2049), .n2048(n2048), 
            .n2047(n2047), .\mem_LUT.mem_3_3 (\mem_LUT.mem_3_3 ), .n2046(n2046), 
            .\mem_LUT.mem_3_2 (\mem_LUT.mem_3_2 ), .n2045(n2045), .\mem_LUT.mem_3_1 (\mem_LUT.mem_3_1 ), 
            .n2044(n2044), .\mem_LUT.mem_3_0 (\mem_LUT.mem_3_0 ), .\mem_LUT.mem_1_6 (\mem_LUT.mem_1_6 ), 
            .n1957(n1957), .\mem_LUT.mem_1_0 (\mem_LUT.mem_1_0 ), .n1954(n1954), 
            .\mem_LUT.mem_1_1 (\mem_LUT.mem_1_1 ), .n1951(n1951), .\mem_LUT.mem_1_2 (\mem_LUT.mem_1_2 ), 
            .n1945(n1945), .\mem_LUT.mem_1_3 (\mem_LUT.mem_1_3 ), .n1944(n1944), 
            .n1939(n1939), .n1935(n1935), .n1930(n1930), .\mem_LUT.mem_1_7 (\mem_LUT.mem_1_7 ), 
            .n1983(n1983), .rd_fifo_en_prev_r(rd_fifo_en_prev_r), .\wr_addr_p1_w[2] (wr_addr_p1_w[2]), 
            .n2968(n2968), .rx_buf_byte({rx_buf_byte}), .RESET_c(RESET_c), 
            .n4(n4_adj_494), .n2(n2), .\rd_addr_p1_w[2] (rd_addr_p1_w[2]), 
            .n3448(n3448), .fifo_read_cmd(fifo_read_cmd)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(604[16] 620[2])
    \uart_tx(CLKS_PER_BIT=434)  pc_tx (.SLM_CLK_c(SLM_CLK_c), .UART_TX_c(UART_TX_c), 
            .r_SM_Main({r_SM_Main_adj_512}), .r_Tx_Data({r_Tx_Data}), .r_Bit_Index({Open_2, 
            Open_3, r_Bit_Index_adj_514[0]}), .GND_net(GND_net), .n3439(n3439), 
            .n2013(n2013), .n2067(n2067), .n2066(n2066), .n2065(n2065), 
            .n2064(n2064), .n2062(n2062), .n2061(n2061), .n2060(n2060), 
            .\r_SM_Main_2__N_187[0] (r_SM_Main_2__N_187[0]), .n1636(n1636), 
            .n1819(n1819), .n1898(n1898), .\r_SM_Main_2__N_184[1] (r_SM_Main_2__N_184[1]), 
            .VCC_net(VCC_net), .n1950(n1950), .n1949(n1949), .tx_uart_active_flag(tx_uart_active_flag), 
            .n4(n4)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(450[42] 459[3])
    
endmodule
//
// Verilog Description of module spi
//

module spi (state_reg, state_next_2__N_312, VCC_net, SDAT_c, reset_all_w, 
            DEBUG_2_c, start_transfer_prev, SLM_CLK_c, n3212, \rx_shift_reg[8] , 
            \tx_shift_reg[0] , n3206, \rx_shift_reg[7] , n3204, \rx_shift_reg[6] , 
            n3198, \rx_shift_reg[5] , SEN_c, n3190, \rx_shift_reg[4] , 
            n3188, \rx_shift_reg[3] , n3184, \rx_shift_reg[2] , n3180, 
            \rx_shift_reg[1] , n2059, \tx_shift_reg[1] , n2057, \tx_shift_reg[2] , 
            n2055, \tx_shift_reg[3] , n2054, \tx_shift_reg[4] , n2053, 
            \tx_shift_reg[5] , n2052, \tx_shift_reg[6] , n2043, \tx_shift_reg[7] , 
            n2042, \tx_shift_reg[8] , n2041, \tx_shift_reg[9] , n2040, 
            \tx_shift_reg[10] , n2039, \tx_shift_reg[11] , n2038, \tx_shift_reg[12] , 
            n2037, \tx_shift_reg[13] , n2036, n2034, rx_buf_byte, 
            n2033, n2032, n2031, n2030, n3148, start_transfer_edge, 
            n2029, n2025, GND_net, spi_busy, n1956, n3178, \rx_shift_reg[0] , 
            n1728, n5, DEBUG_6_c, rx_shift_reg_15__N_319, \tx_data_byte[0] , 
            n883, n3279, \tx_addr_byte[7] ) /* synthesis syn_module_defined=1 */ ;
    output [2:0]state_reg;
    output state_next_2__N_312;
    input VCC_net;
    output SDAT_c;
    input reset_all_w;
    input DEBUG_2_c;
    output start_transfer_prev;
    input SLM_CLK_c;
    input n3212;
    output \rx_shift_reg[8] ;
    output \tx_shift_reg[0] ;
    input n3206;
    output \rx_shift_reg[7] ;
    input n3204;
    output \rx_shift_reg[6] ;
    input n3198;
    output \rx_shift_reg[5] ;
    output SEN_c;
    input n3190;
    output \rx_shift_reg[4] ;
    input n3188;
    output \rx_shift_reg[3] ;
    input n3184;
    output \rx_shift_reg[2] ;
    input n3180;
    output \rx_shift_reg[1] ;
    input n2059;
    output \tx_shift_reg[1] ;
    input n2057;
    output \tx_shift_reg[2] ;
    input n2055;
    output \tx_shift_reg[3] ;
    input n2054;
    output \tx_shift_reg[4] ;
    input n2053;
    output \tx_shift_reg[5] ;
    input n2052;
    output \tx_shift_reg[6] ;
    input n2043;
    output \tx_shift_reg[7] ;
    input n2042;
    output \tx_shift_reg[8] ;
    input n2041;
    output \tx_shift_reg[9] ;
    input n2040;
    output \tx_shift_reg[10] ;
    input n2039;
    output \tx_shift_reg[11] ;
    input n2038;
    output \tx_shift_reg[12] ;
    input n2037;
    output \tx_shift_reg[13] ;
    input n2036;
    input n2034;
    output [7:0]rx_buf_byte;
    input n2033;
    input n2032;
    input n2031;
    input n2030;
    input n3148;
    output start_transfer_edge;
    input n2029;
    input n2025;
    input GND_net;
    output spi_busy;
    input n1956;
    input n3178;
    output \rx_shift_reg[0] ;
    output n1728;
    output n5;
    output DEBUG_6_c;
    output rx_shift_reg_15__N_319;
    input \tx_data_byte[0] ;
    input n883;
    output n3279;
    input \tx_addr_byte[7] ;
    
    wire spi_clk /* synthesis is_clock=1, SET_AS_NETWORK=\spi0/spi_clk */ ;   // src/spi.v(96[5:12])
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n4;
    wire [2:0]state_next;   // src/spi.v(133[10:20])
    wire [15:0]n486;
    wire [15:0]n503;
    
    wire n1731, n3176, spi_clk_N_253, n2431, CS_w, n1679, n890, 
        state_next_2__N_310, state_next_2__N_311;
    wire [15:0]tx_shift_reg;   // src/spi.v(66[26:38])
    
    wire n3328, n906, n1958;
    wire [5:0]n29;
    wire [5:0]spi_clk_counter;   // src/spi.v(97[10:25])
    
    wire n2917, n2919, n2915, n2916, n2918, n1896, n1429, n10, 
        n3337, n2433, n13;
    
    SB_LUT4 i2131_2_lut_4_lut (.I0(state_reg[1]), .I1(n4), .I2(state_next[1]), 
            .I3(n486[4]), .O(n503[5]));   // src/spi.v(165[13:36])
    defparam i2131_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i2130_2_lut_4_lut (.I0(state_reg[1]), .I1(n4), .I2(state_next[1]), 
            .I3(n486[5]), .O(n503[6]));   // src/spi.v(165[13:36])
    defparam i2130_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i2129_2_lut_4_lut (.I0(state_reg[1]), .I1(n4), .I2(state_next[1]), 
            .I3(state_next_2__N_312), .O(n503[7]));   // src/spi.v(165[13:36])
    defparam i2129_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i2128_2_lut_4_lut (.I0(state_reg[1]), .I1(n4), .I2(state_next[1]), 
            .I3(n486[7]), .O(n503[8]));   // src/spi.v(165[13:36])
    defparam i2128_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_DFFNESS tx_shift_reg_i15 (.Q(SDAT_c), .C(spi_clk), .E(VCC_net), 
            .D(n1731), .S(n3176));   // src/spi.v(275[8] 290[4])
    SB_DFFR state_reg_i0 (.Q(state_reg[0]), .C(spi_clk), .D(state_next[0]), 
            .R(reset_all_w));   // src/spi.v(155[10] 157[8])
    SB_DFF start_transfer_prev_74 (.Q(start_transfer_prev), .C(SLM_CLK_c), 
           .D(DEBUG_2_c));   // src/spi.v(73[8] 82[4])
    SB_DFF spi_clk_76 (.Q(spi_clk), .C(SLM_CLK_c), .D(spi_clk_N_253));   // src/spi.v(99[8] 105[44])
    SB_DFF rx__5_i9 (.Q(\rx_shift_reg[8] ), .C(spi_clk), .D(n3212));   // src/spi.v(299[8] 313[4])
    SB_DFFSS CS_w_79 (.Q(CS_w), .C(spi_clk), .D(n2431), .S(state_reg[1]));   // src/spi.v(248[8] 259[4])
    SB_DFFNSR tx_shift_reg_i0 (.Q(\tx_shift_reg[0] ), .C(spi_clk), .D(n1679), 
            .R(n890));   // src/spi.v(275[8] 290[4])
    SB_LUT4 i2127_2_lut_4_lut (.I0(state_reg[1]), .I1(n4), .I2(state_next[1]), 
            .I3(n486[8]), .O(n503[9]));   // src/spi.v(165[13:36])
    defparam i2127_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_DFF rx__5_i8 (.Q(\rx_shift_reg[7] ), .C(spi_clk), .D(n3206));   // src/spi.v(299[8] 313[4])
    SB_DFF rx__5_i7 (.Q(\rx_shift_reg[6] ), .C(spi_clk), .D(n3204));   // src/spi.v(299[8] 313[4])
    SB_DFF rx__5_i6 (.Q(\rx_shift_reg[5] ), .C(spi_clk), .D(n3198));   // src/spi.v(299[8] 313[4])
    SB_DFFS CS_81 (.Q(SEN_c), .C(spi_clk), .D(CS_w), .S(reset_all_w));   // src/spi.v(266[3:14])
    SB_DFFS t_FSM_i0 (.Q(n486[0]), .C(spi_clk), .D(n503[0]), .S(reset_all_w));   // src/spi.v(168[18:23])
    SB_DFF rx__5_i5 (.Q(\rx_shift_reg[4] ), .C(spi_clk), .D(n3190));   // src/spi.v(299[8] 313[4])
    SB_DFF rx__5_i4 (.Q(\rx_shift_reg[3] ), .C(spi_clk), .D(n3188));   // src/spi.v(299[8] 313[4])
    SB_DFF rx__5_i3 (.Q(\rx_shift_reg[2] ), .C(spi_clk), .D(n3184));   // src/spi.v(299[8] 313[4])
    SB_DFF rx__5_i2 (.Q(\rx_shift_reg[1] ), .C(spi_clk), .D(n3180));   // src/spi.v(299[8] 313[4])
    SB_DFFN tx_shift_reg_i1 (.Q(\tx_shift_reg[1] ), .C(spi_clk), .D(n2059));   // src/spi.v(275[8] 290[4])
    SB_DFFN tx_shift_reg_i2 (.Q(\tx_shift_reg[2] ), .C(spi_clk), .D(n2057));   // src/spi.v(275[8] 290[4])
    SB_DFFN tx_shift_reg_i3 (.Q(\tx_shift_reg[3] ), .C(spi_clk), .D(n2055));   // src/spi.v(275[8] 290[4])
    SB_DFFN tx_shift_reg_i4 (.Q(\tx_shift_reg[4] ), .C(spi_clk), .D(n2054));   // src/spi.v(275[8] 290[4])
    SB_DFFN tx_shift_reg_i5 (.Q(\tx_shift_reg[5] ), .C(spi_clk), .D(n2053));   // src/spi.v(275[8] 290[4])
    SB_DFFN tx_shift_reg_i6 (.Q(\tx_shift_reg[6] ), .C(spi_clk), .D(n2052));   // src/spi.v(275[8] 290[4])
    SB_LUT4 i2126_2_lut_4_lut (.I0(state_reg[1]), .I1(n4), .I2(state_next[1]), 
            .I3(n486[9]), .O(n503[10]));   // src/spi.v(165[13:36])
    defparam i2126_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_DFFR t_FSM_i15 (.Q(n486[15]), .C(spi_clk), .D(n503[15]), .R(reset_all_w));   // src/spi.v(168[18:23])
    SB_DFFR t_FSM_i14 (.Q(n486[14]), .C(spi_clk), .D(n503[14]), .R(reset_all_w));   // src/spi.v(168[18:23])
    SB_DFFR t_FSM_i13 (.Q(n486[13]), .C(spi_clk), .D(n503[13]), .R(reset_all_w));   // src/spi.v(168[18:23])
    SB_DFFR t_FSM_i12 (.Q(n486[12]), .C(spi_clk), .D(n503[12]), .R(reset_all_w));   // src/spi.v(168[18:23])
    SB_DFFR t_FSM_i11 (.Q(n486[11]), .C(spi_clk), .D(n503[11]), .R(reset_all_w));   // src/spi.v(168[18:23])
    SB_DFFR t_FSM_i10 (.Q(n486[10]), .C(spi_clk), .D(n503[10]), .R(reset_all_w));   // src/spi.v(168[18:23])
    SB_DFFR t_FSM_i9 (.Q(n486[9]), .C(spi_clk), .D(n503[9]), .R(reset_all_w));   // src/spi.v(168[18:23])
    SB_DFFR t_FSM_i8 (.Q(n486[8]), .C(spi_clk), .D(n503[8]), .R(reset_all_w));   // src/spi.v(168[18:23])
    SB_DFFR t_FSM_i7 (.Q(n486[7]), .C(spi_clk), .D(n503[7]), .R(reset_all_w));   // src/spi.v(168[18:23])
    SB_DFFR t_FSM_i6 (.Q(state_next_2__N_312), .C(spi_clk), .D(n503[6]), 
            .R(reset_all_w));   // src/spi.v(168[18:23])
    SB_DFFR t_FSM_i5 (.Q(n486[5]), .C(spi_clk), .D(n503[5]), .R(reset_all_w));   // src/spi.v(168[18:23])
    SB_DFFR t_FSM_i4 (.Q(n486[4]), .C(spi_clk), .D(n503[4]), .R(reset_all_w));   // src/spi.v(168[18:23])
    SB_DFFN tx_shift_reg_i7 (.Q(\tx_shift_reg[7] ), .C(spi_clk), .D(n2043));   // src/spi.v(275[8] 290[4])
    SB_DFFN tx_shift_reg_i8 (.Q(\tx_shift_reg[8] ), .C(spi_clk), .D(n2042));   // src/spi.v(275[8] 290[4])
    SB_DFFN tx_shift_reg_i9 (.Q(\tx_shift_reg[9] ), .C(spi_clk), .D(n2041));   // src/spi.v(275[8] 290[4])
    SB_DFFN tx_shift_reg_i10 (.Q(\tx_shift_reg[10] ), .C(spi_clk), .D(n2040));   // src/spi.v(275[8] 290[4])
    SB_DFFR t_FSM_i3 (.Q(n486[3]), .C(spi_clk), .D(n503[3]), .R(reset_all_w));   // src/spi.v(168[18:23])
    SB_DFFR t_FSM_i2 (.Q(state_next_2__N_310), .C(spi_clk), .D(n503[2]), 
            .R(reset_all_w));   // src/spi.v(168[18:23])
    SB_DFFR t_FSM_i1 (.Q(state_next_2__N_311), .C(spi_clk), .D(n503[1]), 
            .R(reset_all_w));   // src/spi.v(168[18:23])
    SB_DFFN tx_shift_reg_i11 (.Q(\tx_shift_reg[11] ), .C(spi_clk), .D(n2039));   // src/spi.v(275[8] 290[4])
    SB_DFFN tx_shift_reg_i12 (.Q(\tx_shift_reg[12] ), .C(spi_clk), .D(n2038));   // src/spi.v(275[8] 290[4])
    SB_DFFN tx_shift_reg_i13 (.Q(\tx_shift_reg[13] ), .C(spi_clk), .D(n2037));   // src/spi.v(275[8] 290[4])
    SB_DFFN tx_shift_reg_i14 (.Q(tx_shift_reg[14]), .C(spi_clk), .D(n2036));   // src/spi.v(275[8] 290[4])
    SB_DFF Rx_Lower_Byte_i1 (.Q(rx_buf_byte[1]), .C(spi_clk), .D(n2034));   // src/spi.v(299[8] 313[4])
    SB_DFF Rx_Lower_Byte_i2 (.Q(rx_buf_byte[2]), .C(spi_clk), .D(n2033));   // src/spi.v(299[8] 313[4])
    SB_DFF Rx_Lower_Byte_i3 (.Q(rx_buf_byte[3]), .C(spi_clk), .D(n2032));   // src/spi.v(299[8] 313[4])
    SB_DFF Rx_Lower_Byte_i4 (.Q(rx_buf_byte[4]), .C(spi_clk), .D(n2031));   // src/spi.v(299[8] 313[4])
    SB_DFF Rx_Lower_Byte_i5 (.Q(rx_buf_byte[5]), .C(spi_clk), .D(n2030));   // src/spi.v(299[8] 313[4])
    SB_DFF start_transfer_edge_73 (.Q(start_transfer_edge), .C(SLM_CLK_c), 
           .D(n3148));   // src/spi.v(73[8] 82[4])
    SB_DFFR state_reg_i2 (.Q(state_reg[2]), .C(spi_clk), .D(state_next[2]), 
            .R(reset_all_w));   // src/spi.v(155[10] 157[8])
    SB_DFF Rx_Lower_Byte_i6 (.Q(rx_buf_byte[6]), .C(spi_clk), .D(n2029));   // src/spi.v(299[8] 313[4])
    SB_DFFR state_reg_i1 (.Q(state_reg[1]), .C(spi_clk), .D(state_next[1]), 
            .R(reset_all_w));   // src/spi.v(155[10] 157[8])
    SB_DFF Rx_Lower_Byte_i7 (.Q(rx_buf_byte[7]), .C(spi_clk), .D(n2025));   // src/spi.v(299[8] 313[4])
    SB_LUT4 i2963_2_lut_3_lut (.I0(state_reg[0]), .I1(state_reg[1]), .I2(state_next_2__N_310), 
            .I3(GND_net), .O(n3328));   // src/spi.v(155[10] 157[8])
    defparam i2963_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1_2_lut_3_lut (.I0(state_reg[0]), .I1(state_reg[1]), .I2(state_next_2__N_312), 
            .I3(GND_net), .O(n906));   // src/spi.v(155[10] 157[8])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1_4_lut (.I0(state_reg[2]), .I1(state_reg[0]), .I2(state_next[2]), 
            .I3(state_next[0]), .O(n4));   // src/spi.v(165[13:36])
    defparam i1_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_1_lut (.I0(state_reg[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n890));   // src/spi.v(280[5] 288[12])
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1605_2_lut_3_lut (.I0(state_reg[1]), .I1(state_reg[2]), .I2(state_reg[0]), 
            .I3(GND_net), .O(n1958));   // src/spi.v(282[6:10])
    defparam i1605_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF busy_86 (.Q(spi_busy), .C(spi_clk), .D(n1958));   // src/spi.v(320[8] 326[4])
    SB_LUT4 spi_clk_counter_587_add_4_5_lut (.I0(GND_net), .I1(VCC_net), 
            .I2(spi_clk_counter[3]), .I3(n2917), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam spi_clk_counter_587_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 spi_clk_counter_587_add_4_7_lut (.I0(GND_net), .I1(VCC_net), 
            .I2(spi_clk_counter[5]), .I3(n2919), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam spi_clk_counter_587_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 spi_clk_counter_587_add_4_3_lut (.I0(GND_net), .I1(VCC_net), 
            .I2(spi_clk_counter[1]), .I3(n2915), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam spi_clk_counter_587_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY spi_clk_counter_587_add_4_3 (.CI(n2915), .I0(VCC_net), .I1(spi_clk_counter[1]), 
            .CO(n2916));
    SB_CARRY spi_clk_counter_587_add_4_5 (.CI(n2917), .I0(VCC_net), .I1(spi_clk_counter[3]), 
            .CO(n2918));
    SB_LUT4 spi_clk_counter_587_add_4_4_lut (.I0(GND_net), .I1(VCC_net), 
            .I2(spi_clk_counter[2]), .I3(n2916), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam spi_clk_counter_587_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 spi_clk_counter_587_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(spi_clk_counter[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam spi_clk_counter_587_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR spi_clk_counter_587__i0 (.Q(spi_clk_counter[0]), .C(SLM_CLK_c), 
            .D(n29[0]), .R(n1896));   // src/spi.v(105[21:43])
    SB_LUT4 spi_clk_counter_587_add_4_6_lut (.I0(GND_net), .I1(VCC_net), 
            .I2(spi_clk_counter[4]), .I3(n2918), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam spi_clk_counter_587_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY spi_clk_counter_587_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(spi_clk_counter[0]), 
            .CO(n2915));
    SB_DFF Rx_Lower_Byte_i0 (.Q(rx_buf_byte[0]), .C(spi_clk), .D(n1956));   // src/spi.v(299[8] 313[4])
    SB_DFF rx__5_i1 (.Q(\rx_shift_reg[0] ), .C(spi_clk), .D(n3178));   // src/spi.v(299[8] 313[4])
    SB_DFFSR spi_clk_counter_587__i1 (.Q(spi_clk_counter[1]), .C(SLM_CLK_c), 
            .D(n29[1]), .R(n1896));   // src/spi.v(105[21:43])
    SB_DFFSS spi_clk_counter_587__i2 (.Q(spi_clk_counter[2]), .C(SLM_CLK_c), 
            .D(n29[2]), .S(n1896));   // src/spi.v(105[21:43])
    SB_DFFSR spi_clk_counter_587__i3 (.Q(spi_clk_counter[3]), .C(SLM_CLK_c), 
            .D(n29[3]), .R(n1896));   // src/spi.v(105[21:43])
    SB_DFFSR spi_clk_counter_587__i4 (.Q(spi_clk_counter[4]), .C(SLM_CLK_c), 
            .D(n29[4]), .R(n1896));   // src/spi.v(105[21:43])
    SB_DFFSS spi_clk_counter_587__i5 (.Q(spi_clk_counter[5]), .C(SLM_CLK_c), 
            .D(n29[5]), .S(n1896));   // src/spi.v(105[21:43])
    SB_CARRY spi_clk_counter_587_add_4_4 (.CI(n2916), .I0(VCC_net), .I1(spi_clk_counter[2]), 
            .CO(n2917));
    SB_CARRY spi_clk_counter_587_add_4_6 (.CI(n2918), .I0(VCC_net), .I1(spi_clk_counter[4]), 
            .CO(n2919));
    SB_LUT4 i2125_2_lut_4_lut (.I0(state_reg[1]), .I1(n4), .I2(state_next[1]), 
            .I3(n486[10]), .O(n503[11]));   // src/spi.v(165[13:36])
    defparam i2125_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i1_2_lut_3_lut_adj_14 (.I0(state_reg[0]), .I1(state_reg[2]), 
            .I2(state_reg[1]), .I3(GND_net), .O(n1728));   // src/spi.v(280[5] 288[12])
    defparam i1_2_lut_3_lut_adj_14.LUT_INIT = 16'h0202;
    SB_LUT4 i2_3_lut (.I0(SEN_c), .I1(spi_clk), .I2(n5), .I3(GND_net), 
            .O(DEBUG_6_c));
    defparam i2_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1077_2_lut_4_lut (.I0(state_reg[0]), .I1(state_reg[1]), .I2(state_next_2__N_312), 
            .I3(state_reg[2]), .O(n1429));   // src/spi.v(179[5] 214[12])
    defparam i1077_2_lut_4_lut.LUT_INIT = 16'hdf00;
    SB_LUT4 i2977_2_lut (.I0(state_reg[2]), .I1(state_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n2431));
    defparam i2977_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i2124_2_lut_4_lut (.I0(state_reg[1]), .I1(n4), .I2(state_next[1]), 
            .I3(n486[11]), .O(n503[12]));   // src/spi.v(165[13:36])
    defparam i2124_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i2123_2_lut_4_lut (.I0(state_reg[1]), .I1(n4), .I2(state_next[1]), 
            .I3(n486[12]), .O(n503[13]));   // src/spi.v(165[13:36])
    defparam i2123_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i2122_2_lut_4_lut (.I0(state_reg[1]), .I1(n4), .I2(state_next[1]), 
            .I3(n486[13]), .O(n503[14]));   // src/spi.v(165[13:36])
    defparam i2122_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 state_reg_2__I_0_108_i5_3_lut_3_lut (.I0(state_reg[0]), .I1(state_reg[1]), 
            .I2(state_reg[2]), .I3(GND_net), .O(rx_shift_reg_15__N_319));   // src/spi.v(310[3:14])
    defparam state_reg_2__I_0_108_i5_3_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_15 (.I0(state_reg[2]), .I1(state_reg[1]), 
            .I2(\tx_data_byte[0] ), .I3(GND_net), .O(n1679));   // src/spi.v(280[5] 288[12])
    defparam i1_2_lut_3_lut_adj_15.LUT_INIT = 16'h1010;
    SB_LUT4 i2121_2_lut_4_lut (.I0(state_reg[1]), .I1(n4), .I2(state_next[1]), 
            .I3(n486[14]), .O(n503[15]));   // src/spi.v(165[13:36])
    defparam i2121_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i4_4_lut (.I0(spi_clk_counter[2]), .I1(spi_clk_counter[5]), 
            .I2(spi_clk_counter[0]), .I3(spi_clk_counter[1]), .O(n10));   // src/spi.v(100[5:23])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2987_3_lut (.I0(spi_clk_counter[3]), .I1(n10), .I2(spi_clk_counter[4]), 
            .I3(GND_net), .O(n1896));   // src/spi.v(100[5:23])
    defparam i2987_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_2_lut (.I0(spi_clk), .I1(n1896), .I2(GND_net), .I3(GND_net), 
            .O(spi_clk_N_253));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 state_reg_2__I_0_101_i5_2_lut_3_lut_3_lut (.I0(state_reg[1]), 
            .I1(state_reg[2]), .I2(state_reg[0]), .I3(GND_net), .O(n5));   // src/spi.v(282[6:10])
    defparam state_reg_2__I_0_101_i5_2_lut_3_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i2962_4_lut (.I0(start_transfer_edge), .I1(state_reg[2]), .I2(state_next_2__N_311), 
            .I3(state_reg[1]), .O(n3337));   // src/spi.v(179[5] 214[12])
    defparam i2962_4_lut.LUT_INIT = 16'hcfdd;
    SB_LUT4 i28_4_lut (.I0(n3337), .I1(state_next_2__N_310), .I2(state_reg[0]), 
            .I3(n2433), .O(n13));   // src/spi.v(179[5] 214[12])
    defparam i28_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_512_i1_3_lut (.I0(n13), .I1(n1429), .I2(n883), .I3(GND_net), 
            .O(state_next[0]));   // src/spi.v(179[5] 214[12])
    defparam mux_512_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i2082_2_lut (.I0(state_reg[2]), .I1(state_reg[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2433));
    defparam i2082_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i19_3_lut (.I0(state_reg[1]), .I1(state_reg[2]), .I2(state_reg[0]), 
            .I3(GND_net), .O(n3279));   // src/spi.v(280[5] 288[12])
    defparam i19_3_lut.LUT_INIT = 16'hb9b9;
    SB_LUT4 i1_2_lut_adj_16 (.I0(tx_shift_reg[14]), .I1(n3279), .I2(GND_net), 
            .I3(GND_net), .O(n3176));   // src/spi.v(280[5] 288[12])
    defparam i1_2_lut_adj_16.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_17 (.I0(\tx_addr_byte[7] ), .I1(n1728), .I2(GND_net), 
            .I3(GND_net), .O(n1731));   // src/spi.v(280[5] 288[12])
    defparam i1_2_lut_adj_17.LUT_INIT = 16'h8888;
    SB_LUT4 mux_512_i2_4_lut_4_lut (.I0(state_reg[1]), .I1(state_reg[2]), 
            .I2(n883), .I3(n906), .O(state_next[1]));   // src/spi.v(179[5] 214[12])
    defparam mux_512_i2_4_lut_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 mux_512_i3_4_lut_4_lut (.I0(state_reg[2]), .I1(n883), .I2(n1429), 
            .I3(n3328), .O(state_next[2]));   // src/spi.v(179[5] 214[12])
    defparam mux_512_i3_4_lut_4_lut.LUT_INIT = 16'hf3e2;
    SB_LUT4 i2135_2_lut_4_lut (.I0(state_reg[1]), .I1(n4), .I2(state_next[1]), 
            .I3(n486[0]), .O(n503[1]));   // src/spi.v(165[13:36])
    defparam i2135_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i2134_2_lut_4_lut (.I0(state_reg[1]), .I1(n4), .I2(state_next[1]), 
            .I3(state_next_2__N_311), .O(n503[2]));   // src/spi.v(165[13:36])
    defparam i2134_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i2084_2_lut_4_lut (.I0(state_reg[1]), .I1(n4), .I2(state_next[1]), 
            .I3(n486[15]), .O(n503[0]));   // src/spi.v(165[13:36])
    defparam i2084_2_lut_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i2133_2_lut_4_lut (.I0(state_reg[1]), .I1(n4), .I2(state_next[1]), 
            .I3(state_next_2__N_310), .O(n503[3]));   // src/spi.v(165[13:36])
    defparam i2133_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i2132_2_lut_4_lut (.I0(state_reg[1]), .I1(n4), .I2(state_next[1]), 
            .I3(n486[3]), .O(n503[4]));   // src/spi.v(165[13:36])
    defparam i2132_2_lut_4_lut.LUT_INIT = 16'h2100;
    
endmodule
//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=434) 
//

module \uart_rx(CLKS_PER_BIT=434)  (r_Rx_Data, SLM_CLK_c, n1965, pc_data_rx, 
            \r_SM_Main_2__N_108[2] , GND_net, n3250, r_SM_Main, n2016, 
            r_Bit_Index, n1963, n1962, DEBUG_1_c, n4, n3293, n1747, 
            n2035, uart_rx_complete_prev, n1988, n2540, VCC_net, n1975, 
            n1974, n1973, n1972, UART_RX_c, n1764, n4_adj_3, n1750, 
            n1754, n4_adj_4) /* synthesis syn_module_defined=1 */ ;
    output r_Rx_Data;
    input SLM_CLK_c;
    input n1965;
    output [7:0]pc_data_rx;
    output \r_SM_Main_2__N_108[2] ;
    input GND_net;
    input n3250;
    output [2:0]r_SM_Main;
    input n2016;
    output [2:0]r_Bit_Index;
    input n1963;
    input n1962;
    output DEBUG_1_c;
    output n4;
    output n3293;
    output n1747;
    input n2035;
    input uart_rx_complete_prev;
    output n1988;
    output n2540;
    input VCC_net;
    input n1975;
    input n1974;
    input n1973;
    input n1972;
    input UART_RX_c;
    input n1764;
    output n4_adj_3;
    output n1750;
    output n1754;
    output n4_adj_4;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire r_Rx_Data_R;
    wire [9:0]n45;
    
    wire n1815;
    wire [9:0]r_Clock_Count;   // src/uart_rx.v(32[17:30])
    
    wire n1910, n3261, n2558, n3260, n6, n3291;
    wire [2:0]r_SM_Main_2__N_114;
    
    wire n3271, n3028;
    wire [2:0]r_Bit_Index_c;   // src/uart_rx.v(33[17:28])
    wire [2:0]n340;
    
    wire n1900, n1715, n3334, n3273, n2586, n3, n2922, n2923, 
        n2920, n2921, n2928, n2927, n2926, n2925, n2924, n2578, 
        n1, n6_adj_492;
    
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(SLM_CLK_c), .D(r_Rx_Data_R));   // src/uart_rx.v(41[10] 45[8])
    SB_DFFESR r_Clock_Count_584__i3 (.Q(r_Clock_Count[3]), .C(SLM_CLK_c), 
            .E(n1815), .D(n45[3]), .R(n1910));   // src/uart_rx.v(120[34:51])
    SB_DFF r_Rx_Byte_i3 (.Q(pc_data_rx[3]), .C(SLM_CLK_c), .D(n1965));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_584__i9 (.Q(r_Clock_Count[9]), .C(SLM_CLK_c), 
            .E(n1815), .D(n45[9]), .R(n1910));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_584__i2 (.Q(r_Clock_Count[2]), .C(SLM_CLK_c), 
            .E(n1815), .D(n45[2]), .R(n1910));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_584__i8 (.Q(r_Clock_Count[8]), .C(SLM_CLK_c), 
            .E(n1815), .D(n45[8]), .R(n1910));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_584__i1 (.Q(r_Clock_Count[1]), .C(SLM_CLK_c), 
            .E(n1815), .D(n45[1]), .R(n1910));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_584__i7 (.Q(r_Clock_Count[7]), .C(SLM_CLK_c), 
            .E(n1815), .D(n45[7]), .R(n1910));   // src/uart_rx.v(120[34:51])
    SB_LUT4 i2206_4_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[6]), .I2(n3261), 
            .I3(r_Clock_Count[4]), .O(n2558));
    defparam i2206_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i2220_4_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[9]), .I2(n2558), 
            .I3(r_Clock_Count[7]), .O(\r_SM_Main_2__N_108[2] ));
    defparam i2220_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1_3_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[1]), 
            .I3(GND_net), .O(n3260));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2904_4_lut (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[6]), .I2(r_Clock_Count[3]), 
            .I3(r_Clock_Count[4]), .O(n3291));
    defparam i2904_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[9]), .I1(n3260), .I2(n3291), .I3(n6), 
            .O(r_SM_Main_2__N_114[0]));
    defparam i4_4_lut.LUT_INIT = 16'hffef;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(SLM_CLK_c), .D(n3250));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(SLM_CLK_c), .D(n2016));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2885_2_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_114[0]), .I2(GND_net), 
            .I3(GND_net), .O(n3271));
    defparam i2885_2_lut.LUT_INIT = 16'heeee;
    SB_DFF r_Rx_Byte_i2 (.Q(pc_data_rx[2]), .C(SLM_CLK_c), .D(n1963));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(pc_data_rx[1]), .C(SLM_CLK_c), .D(n1962));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(DEBUG_1_c), .C(SLM_CLK_c), .D(n3028));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 equal_257_i4_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // src/uart_rx.v(97[17:39])
    defparam equal_257_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index_c[1]), .C(SLM_CLK_c), .E(n3293), 
            .D(n340[1]), .R(n1900));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index_c[2]), .C(SLM_CLK_c), .E(n3293), 
            .D(n340[2]), .R(n1900));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index_c[2]), .I1(n1715), .I2(r_Bit_Index_c[1]), 
            .I3(GND_net), .O(n1747));
    defparam i2_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(n3334), 
            .I3(r_SM_Main[1]), .O(n1900));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_4_lut.LUT_INIT = 16'h5011;
    SB_LUT4 i1_4_lut_adj_10 (.I0(r_SM_Main[2]), .I1(n3273), .I2(\r_SM_Main_2__N_108[2] ), 
            .I3(r_SM_Main[1]), .O(n1910));
    defparam i1_4_lut_adj_10.LUT_INIT = 16'h5011;
    SB_DFFESR r_Clock_Count_584__i6 (.Q(r_Clock_Count[6]), .C(SLM_CLK_c), 
            .E(n1815), .D(n45[6]), .R(n1910));   // src/uart_rx.v(120[34:51])
    SB_DFF r_Rx_Byte_i0 (.Q(pc_data_rx[0]), .C(SLM_CLK_c), .D(n2035));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1_2_lut_adj_11 (.I0(DEBUG_1_c), .I1(uart_rx_complete_prev), 
            .I2(GND_net), .I3(GND_net), .O(n1988));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_adj_11.LUT_INIT = 16'h2222;
    SB_LUT4 i706_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n340[1]));   // src/uart_rx.v(102[36:51])
    defparam i706_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2957_2_lut_3_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_108[2] ), 
            .I2(n2540), .I3(GND_net), .O(n3334));   // src/uart_rx.v(52[7] 143[14])
    defparam i2957_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_DFFESR r_Clock_Count_584__i5 (.Q(r_Clock_Count[5]), .C(SLM_CLK_c), 
            .E(n1815), .D(n45[5]), .R(n1910));   // src/uart_rx.v(120[34:51])
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_108[2] ), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[1]), .O(n1715));   // src/uart_rx.v(52[7] 143[14])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_DFFESR r_Clock_Count_584__i4 (.Q(r_Clock_Count[4]), .C(SLM_CLK_c), 
            .E(n1815), .D(n45[4]), .R(n1910));   // src/uart_rx.v(120[34:51])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(SLM_CLK_c), .D(n2586), 
            .R(r_SM_Main[2]));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(SLM_CLK_c), .D(n3), .R(r_SM_Main[2]));   // src/uart_rx.v(49[10] 144[8])
    SB_CARRY r_Clock_Count_584_add_4_5 (.CI(n2922), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n2923));
    SB_CARRY r_Clock_Count_584_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n2920));
    SB_LUT4 r_Clock_Count_584_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[2]), 
            .I3(n2921), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_584_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_584_add_4_4 (.CI(n2921), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n2922));
    SB_LUT4 r_Clock_Count_584_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[1]), 
            .I3(n2920), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_584_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_584_add_4_3 (.CI(n2920), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n2921));
    SB_LUT4 r_Clock_Count_584_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_584_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_584_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[9]), .I3(n2928), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_584_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_584_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n2927), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_584_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_584_add_4_10 (.CI(n2927), .I0(GND_net), .I1(r_Clock_Count[8]), 
            .CO(n2928));
    SB_LUT4 r_Clock_Count_584_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[7]), 
            .I3(n2926), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_584_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_584_add_4_9 (.CI(n2926), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n2927));
    SB_LUT4 r_Clock_Count_584_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[6]), 
            .I3(n2925), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_584_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_584_add_4_8 (.CI(n2925), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n2926));
    SB_LUT4 r_Clock_Count_584_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[5]), 
            .I3(n2924), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_584_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Clock_Count_584__i0 (.Q(r_Clock_Count[0]), .C(SLM_CLK_c), 
            .E(n1815), .D(n45[0]), .R(n1910));   // src/uart_rx.v(120[34:51])
    SB_DFF r_Rx_Byte_i7 (.Q(pc_data_rx[7]), .C(SLM_CLK_c), .D(n1975));   // src/uart_rx.v(49[10] 144[8])
    SB_CARRY r_Clock_Count_584_add_4_7 (.CI(n2924), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n2925));
    SB_DFF r_Rx_Byte_i6 (.Q(pc_data_rx[6]), .C(SLM_CLK_c), .D(n1974));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(pc_data_rx[5]), .C(SLM_CLK_c), .D(n1973));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_Clock_Count_584_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[4]), 
            .I3(n2923), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_584_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i4 (.Q(pc_data_rx[4]), .C(SLM_CLK_c), .D(n1972));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(SLM_CLK_c), .D(UART_RX_c));   // src/uart_rx.v(41[10] 45[8])
    SB_CARRY r_Clock_Count_584_add_4_6 (.CI(n2923), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n2924));
    SB_LUT4 r_Clock_Count_584_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[3]), 
            .I3(n2922), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_584_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_4_lut (.I0(DEBUG_1_c), .I1(r_SM_Main[2]), .I2(n1764), 
            .I3(r_SM_Main[1]), .O(n3028));   // src/uart_rx.v(36[17:26])
    defparam i13_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 equal_261_i4_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_3));   // src/uart_rx.v(97[17:39])
    defparam equal_261_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_12 (.I0(r_Bit_Index[0]), .I1(n1715), .I2(GND_net), 
            .I3(GND_net), .O(n1750));
    defparam i1_2_lut_adj_12.LUT_INIT = 16'heeee;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n2540), .I1(\r_SM_Main_2__N_108[2] ), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n2578));   // src/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_114[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // src/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i3_3_lut (.I0(n1), .I1(n2578), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // src/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_108[2] ), 
            .I2(r_SM_Main[1]), .I3(n3271), .O(n2586));   // src/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h707a;
    SB_LUT4 i2_2_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_114[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_492));
    defparam i2_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2981_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6_adj_492), 
            .I3(r_SM_Main[0]), .O(n1815));   // src/uart_rx.v(52[7] 143[14])
    defparam i2981_4_lut.LUT_INIT = 16'h4555;
    SB_LUT4 i713_2_lut_3_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), 
            .I2(r_Bit_Index_c[2]), .I3(GND_net), .O(n340[2]));   // src/uart_rx.v(102[36:51])
    defparam i713_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), 
            .I2(r_Bit_Index_c[2]), .I3(GND_net), .O(n2540));   // src/uart_rx.v(102[36:51])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2996_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_108[2] ), .O(n3293));
    defparam i2996_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i2887_2_lut_3_lut (.I0(r_SM_Main[0]), .I1(r_Rx_Data), .I2(r_SM_Main_2__N_114[0]), 
            .I3(GND_net), .O(n3273));
    defparam i2887_2_lut_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_2_lut_4_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[0]), 
            .I2(r_Clock_Count[2]), .I3(r_Clock_Count[1]), .O(n3261));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_13 (.I0(n1715), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1754));   // src/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_13.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_258_i4_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4));   // src/uart_rx.v(97[17:39])
    defparam equal_258_i4_2_lut.LUT_INIT = 16'hdddd;
    
endmodule
//
// Verilog Description of module clock
//

module clock (GND_net, VCC_net, ICE_SYSCLK_c, pll_clk_unbuf) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    input ICE_SYSCLK_c;
    output pll_clk_unbuf;
    
    
    SB_PLL40_CORE pll_config (.REFERENCECLK(ICE_SYSCLK_c), .PLLOUTGLOBAL(pll_clk_unbuf), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=214, LSE_RLINE=219 */ ;   // src/top.v(214[7] 219[3])
    defparam pll_config.FEEDBACK_PATH = "SIMPLE";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll_config.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll_config.FDA_FEEDBACK = 0;
    defparam pll_config.FDA_RELATIVE = 0;
    defparam pll_config.PLLOUT_SELECT = "GENCLK";
    defparam pll_config.DIVR = 4'b0001;
    defparam pll_config.DIVF = 7'b1000010;
    defparam pll_config.DIVQ = 3'b100;
    defparam pll_config.FILTER_RANGE = 3'b001;
    defparam pll_config.ENABLE_ICEGATE = 1'b0;
    defparam pll_config.TEST_MODE = 1'b0;
    defparam pll_config.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module FIFO_Quad_Word
//

module FIFO_Quad_Word (rd_fifo_en_w, \mem_LUT.data_raw_r[0] , SLM_CLK_c, 
            n3239, is_fifo_empty_flag, n1968, \fifo_temp_output[5] , 
            rd_addr_r, \mem_LUT.mem_3_5 , n1971, \fifo_temp_output[6] , 
            \mem_LUT.mem_1_5 , n1978, n1981, n3118, is_tx_fifo_full_flag, 
            n1933, \fifo_temp_output[3] , n1994, \fifo_temp_output[7] , 
            n1938, wr_addr_r, n1942, \fifo_temp_output[4] , n8, reset_all_w, 
            n1948, n8_adj_2, n2009, \fifo_temp_output[0] , fifo_write_cmd, 
            wr_fifo_en_w, GND_net, n2076, VCC_net, \fifo_temp_output[2] , 
            n2073, \fifo_temp_output[1] , \mem_LUT.data_raw_r[7] , n1, 
            \mem_LUT.data_raw_r[6] , \mem_LUT.data_raw_r[5] , \mem_LUT.data_raw_r[4] , 
            \mem_LUT.data_raw_r[3] , \mem_LUT.data_raw_r[2] , \mem_LUT.data_raw_r[1] , 
            n2051, \mem_LUT.mem_3_7 , n2050, \mem_LUT.mem_3_6 , \mem_LUT.mem_3_4 , 
            \mem_LUT.mem_1_4 , n2049, n2048, n2047, \mem_LUT.mem_3_3 , 
            n2046, \mem_LUT.mem_3_2 , n2045, \mem_LUT.mem_3_1 , n2044, 
            \mem_LUT.mem_3_0 , \mem_LUT.mem_1_6 , n1957, \mem_LUT.mem_1_0 , 
            n1954, \mem_LUT.mem_1_1 , n1951, \mem_LUT.mem_1_2 , n1945, 
            \mem_LUT.mem_1_3 , n1944, n1939, n1935, n1930, \mem_LUT.mem_1_7 , 
            n1983, rd_fifo_en_prev_r, \wr_addr_p1_w[2] , n2968, rx_buf_byte, 
            RESET_c, n4, n2, \rd_addr_p1_w[2] , n3448, fifo_read_cmd) /* synthesis syn_module_defined=1 */ ;
    output rd_fifo_en_w;
    output \mem_LUT.data_raw_r[0] ;
    input SLM_CLK_c;
    input n3239;
    output is_fifo_empty_flag;
    input n1968;
    output \fifo_temp_output[5] ;
    output [2:0]rd_addr_r;
    output \mem_LUT.mem_3_5 ;
    input n1971;
    output \fifo_temp_output[6] ;
    output \mem_LUT.mem_1_5 ;
    input n1978;
    input n1981;
    input n3118;
    output is_tx_fifo_full_flag;
    input n1933;
    output \fifo_temp_output[3] ;
    input n1994;
    output \fifo_temp_output[7] ;
    input n1938;
    output [2:0]wr_addr_r;
    input n1942;
    output \fifo_temp_output[4] ;
    input n8;
    input reset_all_w;
    input n1948;
    input n8_adj_2;
    input n2009;
    output \fifo_temp_output[0] ;
    input fifo_write_cmd;
    output wr_fifo_en_w;
    input GND_net;
    input n2076;
    input VCC_net;
    output \fifo_temp_output[2] ;
    input n2073;
    output \fifo_temp_output[1] ;
    output \mem_LUT.data_raw_r[7] ;
    output n1;
    output \mem_LUT.data_raw_r[6] ;
    output \mem_LUT.data_raw_r[5] ;
    output \mem_LUT.data_raw_r[4] ;
    output \mem_LUT.data_raw_r[3] ;
    output \mem_LUT.data_raw_r[2] ;
    output \mem_LUT.data_raw_r[1] ;
    input n2051;
    output \mem_LUT.mem_3_7 ;
    input n2050;
    output \mem_LUT.mem_3_6 ;
    output \mem_LUT.mem_3_4 ;
    output \mem_LUT.mem_1_4 ;
    input n2049;
    input n2048;
    input n2047;
    output \mem_LUT.mem_3_3 ;
    input n2046;
    output \mem_LUT.mem_3_2 ;
    input n2045;
    output \mem_LUT.mem_3_1 ;
    input n2044;
    output \mem_LUT.mem_3_0 ;
    output \mem_LUT.mem_1_6 ;
    input n1957;
    output \mem_LUT.mem_1_0 ;
    input n1954;
    output \mem_LUT.mem_1_1 ;
    input n1951;
    output \mem_LUT.mem_1_2 ;
    input n1945;
    output \mem_LUT.mem_1_3 ;
    input n1944;
    input n1939;
    input n1935;
    input n1930;
    output \mem_LUT.mem_1_7 ;
    input n1983;
    output rd_fifo_en_prev_r;
    output \wr_addr_p1_w[2] ;
    output n2968;
    input [7:0]rx_buf_byte;
    output RESET_c;
    output n4;
    output n2;
    output \rd_addr_p1_w[2] ;
    output n3448;
    input fifo_read_cmd;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_1 lscc_fifo_inst (.rd_fifo_en_w(rd_fifo_en_w), 
            .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r[0] ), .SLM_CLK_c(SLM_CLK_c), 
            .n3239(n3239), .is_fifo_empty_flag(is_fifo_empty_flag), .n1968(n1968), 
            .\fifo_temp_output[5] (\fifo_temp_output[5] ), .rd_addr_r({rd_addr_r}), 
            .\mem_LUT.mem_3_5 (\mem_LUT.mem_3_5 ), .n1971(n1971), .\fifo_temp_output[6] (\fifo_temp_output[6] ), 
            .\mem_LUT.mem_1_5 (\mem_LUT.mem_1_5 ), .n1978(n1978), .n1981(n1981), 
            .n3118(n3118), .is_tx_fifo_full_flag(is_tx_fifo_full_flag), 
            .n1933(n1933), .\fifo_temp_output[3] (\fifo_temp_output[3] ), 
            .n1994(n1994), .\fifo_temp_output[7] (\fifo_temp_output[7] ), 
            .n1938(n1938), .wr_addr_r({wr_addr_r}), .n1942(n1942), .\fifo_temp_output[4] (\fifo_temp_output[4] ), 
            .n8(n8), .reset_all_w(reset_all_w), .n1948(n1948), .n8_adj_1(n8_adj_2), 
            .n2009(n2009), .\fifo_temp_output[0] (\fifo_temp_output[0] ), 
            .fifo_write_cmd(fifo_write_cmd), .wr_fifo_en_w(wr_fifo_en_w), 
            .GND_net(GND_net), .n2076(n2076), .VCC_net(VCC_net), .\fifo_temp_output[2] (\fifo_temp_output[2] ), 
            .n2073(n2073), .\fifo_temp_output[1] (\fifo_temp_output[1] ), 
            .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r[7] ), .n1(n1), 
            .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r[6] ), .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r[5] ), 
            .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r[4] ), .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r[3] ), 
            .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r[2] ), .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r[1] ), 
            .n2051(n2051), .\mem_LUT.mem_3_7 (\mem_LUT.mem_3_7 ), .n2050(n2050), 
            .\mem_LUT.mem_3_6 (\mem_LUT.mem_3_6 ), .\mem_LUT.mem_3_4 (\mem_LUT.mem_3_4 ), 
            .\mem_LUT.mem_1_4 (\mem_LUT.mem_1_4 ), .n2049(n2049), .n2048(n2048), 
            .n2047(n2047), .\mem_LUT.mem_3_3 (\mem_LUT.mem_3_3 ), .n2046(n2046), 
            .\mem_LUT.mem_3_2 (\mem_LUT.mem_3_2 ), .n2045(n2045), .\mem_LUT.mem_3_1 (\mem_LUT.mem_3_1 ), 
            .n2044(n2044), .\mem_LUT.mem_3_0 (\mem_LUT.mem_3_0 ), .\mem_LUT.mem_1_6 (\mem_LUT.mem_1_6 ), 
            .n1957(n1957), .\mem_LUT.mem_1_0 (\mem_LUT.mem_1_0 ), .n1954(n1954), 
            .\mem_LUT.mem_1_1 (\mem_LUT.mem_1_1 ), .n1951(n1951), .\mem_LUT.mem_1_2 (\mem_LUT.mem_1_2 ), 
            .n1945(n1945), .\mem_LUT.mem_1_3 (\mem_LUT.mem_1_3 ), .n1944(n1944), 
            .n1939(n1939), .n1935(n1935), .n1930(n1930), .\mem_LUT.mem_1_7 (\mem_LUT.mem_1_7 ), 
            .n1983(n1983), .rd_fifo_en_prev_r(rd_fifo_en_prev_r), .\wr_addr_p1_w[2] (\wr_addr_p1_w[2] ), 
            .n2968(n2968), .rx_buf_byte({rx_buf_byte}), .RESET_c(RESET_c), 
            .n4(n4), .n2(n2), .\rd_addr_p1_w[2] (\rd_addr_p1_w[2] ), .n3448(n3448), 
            .fifo_read_cmd(fifo_read_cmd)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_quad_word_mod.v(20[37:380])
    
endmodule
//
// Verilog Description of module FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_1
//

module FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_1 (rd_fifo_en_w, 
            \mem_LUT.data_raw_r[0] , SLM_CLK_c, n3239, is_fifo_empty_flag, 
            n1968, \fifo_temp_output[5] , rd_addr_r, \mem_LUT.mem_3_5 , 
            n1971, \fifo_temp_output[6] , \mem_LUT.mem_1_5 , n1978, 
            n1981, n3118, is_tx_fifo_full_flag, n1933, \fifo_temp_output[3] , 
            n1994, \fifo_temp_output[7] , n1938, wr_addr_r, n1942, 
            \fifo_temp_output[4] , n8, reset_all_w, n1948, n8_adj_1, 
            n2009, \fifo_temp_output[0] , fifo_write_cmd, wr_fifo_en_w, 
            GND_net, n2076, VCC_net, \fifo_temp_output[2] , n2073, 
            \fifo_temp_output[1] , \mem_LUT.data_raw_r[7] , n1, \mem_LUT.data_raw_r[6] , 
            \mem_LUT.data_raw_r[5] , \mem_LUT.data_raw_r[4] , \mem_LUT.data_raw_r[3] , 
            \mem_LUT.data_raw_r[2] , \mem_LUT.data_raw_r[1] , n2051, \mem_LUT.mem_3_7 , 
            n2050, \mem_LUT.mem_3_6 , \mem_LUT.mem_3_4 , \mem_LUT.mem_1_4 , 
            n2049, n2048, n2047, \mem_LUT.mem_3_3 , n2046, \mem_LUT.mem_3_2 , 
            n2045, \mem_LUT.mem_3_1 , n2044, \mem_LUT.mem_3_0 , \mem_LUT.mem_1_6 , 
            n1957, \mem_LUT.mem_1_0 , n1954, \mem_LUT.mem_1_1 , n1951, 
            \mem_LUT.mem_1_2 , n1945, \mem_LUT.mem_1_3 , n1944, n1939, 
            n1935, n1930, \mem_LUT.mem_1_7 , n1983, rd_fifo_en_prev_r, 
            \wr_addr_p1_w[2] , n2968, rx_buf_byte, RESET_c, n4, n2, 
            \rd_addr_p1_w[2] , n3448, fifo_read_cmd) /* synthesis syn_module_defined=1 */ ;
    output rd_fifo_en_w;
    output \mem_LUT.data_raw_r[0] ;
    input SLM_CLK_c;
    input n3239;
    output is_fifo_empty_flag;
    input n1968;
    output \fifo_temp_output[5] ;
    output [2:0]rd_addr_r;
    output \mem_LUT.mem_3_5 ;
    input n1971;
    output \fifo_temp_output[6] ;
    output \mem_LUT.mem_1_5 ;
    input n1978;
    input n1981;
    input n3118;
    output is_tx_fifo_full_flag;
    input n1933;
    output \fifo_temp_output[3] ;
    input n1994;
    output \fifo_temp_output[7] ;
    input n1938;
    output [2:0]wr_addr_r;
    input n1942;
    output \fifo_temp_output[4] ;
    input n8;
    input reset_all_w;
    input n1948;
    input n8_adj_1;
    input n2009;
    output \fifo_temp_output[0] ;
    input fifo_write_cmd;
    output wr_fifo_en_w;
    input GND_net;
    input n2076;
    input VCC_net;
    output \fifo_temp_output[2] ;
    input n2073;
    output \fifo_temp_output[1] ;
    output \mem_LUT.data_raw_r[7] ;
    output n1;
    output \mem_LUT.data_raw_r[6] ;
    output \mem_LUT.data_raw_r[5] ;
    output \mem_LUT.data_raw_r[4] ;
    output \mem_LUT.data_raw_r[3] ;
    output \mem_LUT.data_raw_r[2] ;
    output \mem_LUT.data_raw_r[1] ;
    input n2051;
    output \mem_LUT.mem_3_7 ;
    input n2050;
    output \mem_LUT.mem_3_6 ;
    output \mem_LUT.mem_3_4 ;
    output \mem_LUT.mem_1_4 ;
    input n2049;
    input n2048;
    input n2047;
    output \mem_LUT.mem_3_3 ;
    input n2046;
    output \mem_LUT.mem_3_2 ;
    input n2045;
    output \mem_LUT.mem_3_1 ;
    input n2044;
    output \mem_LUT.mem_3_0 ;
    output \mem_LUT.mem_1_6 ;
    input n1957;
    output \mem_LUT.mem_1_0 ;
    input n1954;
    output \mem_LUT.mem_1_1 ;
    input n1951;
    output \mem_LUT.mem_1_2 ;
    input n1945;
    output \mem_LUT.mem_1_3 ;
    input n1944;
    input n1939;
    input n1935;
    input n1930;
    output \mem_LUT.mem_1_7 ;
    input n1983;
    output rd_fifo_en_prev_r;
    output \wr_addr_p1_w[2] ;
    output n2968;
    input [7:0]rx_buf_byte;
    output RESET_c;
    output n4;
    output n2;
    output \rd_addr_p1_w[2] ;
    output n3448;
    input fifo_read_cmd;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [31:0]\mem_LUT.data_raw_r_31__N_402 ;
    
    wire \mem_LUT.mem_2_5 , n3409, \mem_LUT.mem_0_5 , \mem_LUT.mem_2_4 , 
        n3403, \mem_LUT.mem_0_4 , \mem_LUT.mem_2_6 , n3397, n1959, 
        \mem_LUT.mem_0_0 , \mem_LUT.mem_0_6 , n2024, \mem_LUT.mem_2_7 , 
        n2023, n2022, n2021, n2020, \mem_LUT.mem_2_3 , n2019, \mem_LUT.mem_2_2 , 
        n2018, \mem_LUT.mem_2_1 , n2017, \mem_LUT.mem_2_0 , n1955, 
        \mem_LUT.mem_0_1 , n1953, \mem_LUT.mem_0_2 , n1952, \mem_LUT.mem_0_3 , 
        n3391, n1943, n1934, n1928, \mem_LUT.mem_0_7 , n1927, n2_c, 
        n4_c, n3433, n3427, n3421, n3415;
    
    SB_DFFE \mem_LUT.data_raw_r__i1  (.Q(\mem_LUT.data_raw_r[0] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_402 [0]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFF empty_r_85 (.Q(is_fifo_empty_flag), .C(SLM_CLK_c), .D(n3239));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF \mem_LUT.data_buff_r__i5  (.Q(\fifo_temp_output[5] ), .C(SLM_CLK_c), 
           .D(n1968));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_3024 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_5 ), 
            .I2(\mem_LUT.mem_3_5 ), .I3(rd_addr_r[1]), .O(n3409));
    defparam rd_addr_r_0__bdd_4_lut_3024.LUT_INIT = 16'he4aa;
    SB_DFF \mem_LUT.data_buff_r__i6  (.Q(\fifo_temp_output[6] ), .C(SLM_CLK_c), 
           .D(n1971));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 n3409_bdd_4_lut (.I0(n3409), .I1(\mem_LUT.mem_1_5 ), .I2(\mem_LUT.mem_0_5 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_402 [5]));
    defparam n3409_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF rd_addr_r__i1 (.Q(rd_addr_r[1]), .C(SLM_CLK_c), .D(n1978));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF rd_addr_r__i2 (.Q(rd_addr_r[2]), .C(SLM_CLK_c), .D(n1981));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF full_r_84 (.Q(is_tx_fifo_full_flag), .C(SLM_CLK_c), .D(n3118));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF \mem_LUT.data_buff_r__i3  (.Q(\fifo_temp_output[3] ), .C(SLM_CLK_c), 
           .D(n1933));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i7  (.Q(\fifo_temp_output[7] ), .C(SLM_CLK_c), 
           .D(n1994));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF wr_addr_r__i1 (.Q(wr_addr_r[1]), .C(SLM_CLK_c), .D(n1938));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF \mem_LUT.data_buff_r__i4  (.Q(\fifo_temp_output[4] ), .C(SLM_CLK_c), 
           .D(n1942));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFSR wr_addr_r__i0 (.Q(wr_addr_r[0]), .C(SLM_CLK_c), .D(n8), .R(reset_all_w));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF wr_addr_r__i2 (.Q(wr_addr_r[2]), .C(SLM_CLK_c), .D(n1948));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFSR rd_addr_r__i0 (.Q(rd_addr_r[0]), .C(SLM_CLK_c), .D(n8_adj_1), 
            .R(reset_all_w));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF \mem_LUT.data_buff_r__i0  (.Q(\fifo_temp_output[0] ), .C(SLM_CLK_c), 
           .D(n2009));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 wr_en_i_I_0_2_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(GND_net), .I3(GND_net), .O(wr_fifo_en_w));   // src/fifo_quad_word_mod.v(103[21:60])
    defparam wr_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE \mem_LUT.data_buff_r__i2  (.Q(\fifo_temp_output[2] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n2076));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE \mem_LUT.data_buff_r__i1  (.Q(\fifo_temp_output[1] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n2073));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE \mem_LUT.data_raw_r__i8  (.Q(\mem_LUT.data_raw_r[7] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_402 [7]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_LUT4 wr_addr_r_1__I_0_i1_2_lut (.I0(wr_addr_r[0]), .I1(rd_addr_r[0]), 
            .I2(GND_net), .I3(GND_net), .O(n1));   // src/fifo_quad_word_mod.v(115[26:58])
    defparam wr_addr_r_1__I_0_i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE \mem_LUT.data_raw_r__i7  (.Q(\mem_LUT.data_raw_r[6] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_402 [6]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i6  (.Q(\mem_LUT.data_raw_r[5] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_402 [5]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i5  (.Q(\mem_LUT.data_raw_r[4] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_402 [4]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i4  (.Q(\mem_LUT.data_raw_r[3] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_402 [3]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i3  (.Q(\mem_LUT.data_raw_r[2] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_402 [2]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i2  (.Q(\mem_LUT.data_raw_r[1] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_402 [1]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFF i347_348 (.Q(\mem_LUT.mem_3_7 ), .C(SLM_CLK_c), .D(n2051));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i344_345 (.Q(\mem_LUT.mem_3_6 ), .C(SLM_CLK_c), .D(n2050));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_3019 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_4 ), 
            .I2(\mem_LUT.mem_3_4 ), .I3(rd_addr_r[1]), .O(n3403));
    defparam rd_addr_r_0__bdd_4_lut_3019.LUT_INIT = 16'he4aa;
    SB_LUT4 n3403_bdd_4_lut (.I0(n3403), .I1(\mem_LUT.mem_1_4 ), .I2(\mem_LUT.mem_0_4 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_402 [4]));
    defparam n3403_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i341_342 (.Q(\mem_LUT.mem_3_5 ), .C(SLM_CLK_c), .D(n2049));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i338_339 (.Q(\mem_LUT.mem_3_4 ), .C(SLM_CLK_c), .D(n2048));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i335_336 (.Q(\mem_LUT.mem_3_3 ), .C(SLM_CLK_c), .D(n2047));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i332_333 (.Q(\mem_LUT.mem_3_2 ), .C(SLM_CLK_c), .D(n2046));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i329_330 (.Q(\mem_LUT.mem_3_1 ), .C(SLM_CLK_c), .D(n2045));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i326_327 (.Q(\mem_LUT.mem_3_0 ), .C(SLM_CLK_c), .D(n2044));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_3014 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_6 ), 
            .I2(\mem_LUT.mem_3_6 ), .I3(rd_addr_r[1]), .O(n3397));
    defparam rd_addr_r_0__bdd_4_lut_3014.LUT_INIT = 16'he4aa;
    SB_DFF i38_39 (.Q(\mem_LUT.mem_0_0 ), .C(SLM_CLK_c), .D(n1959));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 n3397_bdd_4_lut (.I0(n3397), .I1(\mem_LUT.mem_1_6 ), .I2(\mem_LUT.mem_0_6 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_402 [6]));
    defparam n3397_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i251_252 (.Q(\mem_LUT.mem_2_7 ), .C(SLM_CLK_c), .D(n2024));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i248_249 (.Q(\mem_LUT.mem_2_6 ), .C(SLM_CLK_c), .D(n2023));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i245_246 (.Q(\mem_LUT.mem_2_5 ), .C(SLM_CLK_c), .D(n2022));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i242_243 (.Q(\mem_LUT.mem_2_4 ), .C(SLM_CLK_c), .D(n2021));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i239_240 (.Q(\mem_LUT.mem_2_3 ), .C(SLM_CLK_c), .D(n2020));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i236_237 (.Q(\mem_LUT.mem_2_2 ), .C(SLM_CLK_c), .D(n2019));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i233_234 (.Q(\mem_LUT.mem_2_1 ), .C(SLM_CLK_c), .D(n2018));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i230_231 (.Q(\mem_LUT.mem_2_0 ), .C(SLM_CLK_c), .D(n2017));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i134_135 (.Q(\mem_LUT.mem_1_0 ), .C(SLM_CLK_c), .D(n1957));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i41_42 (.Q(\mem_LUT.mem_0_1 ), .C(SLM_CLK_c), .D(n1955));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i137_138 (.Q(\mem_LUT.mem_1_1 ), .C(SLM_CLK_c), .D(n1954));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i44_45 (.Q(\mem_LUT.mem_0_2 ), .C(SLM_CLK_c), .D(n1953));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i47_48 (.Q(\mem_LUT.mem_0_3 ), .C(SLM_CLK_c), .D(n1952));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i140_141 (.Q(\mem_LUT.mem_1_2 ), .C(SLM_CLK_c), .D(n1951));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i143_144 (.Q(\mem_LUT.mem_1_3 ), .C(SLM_CLK_c), .D(n1945));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i146_147 (.Q(\mem_LUT.mem_1_4 ), .C(SLM_CLK_c), .D(n1944));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_3009 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_3 ), 
            .I2(\mem_LUT.mem_3_3 ), .I3(rd_addr_r[1]), .O(n3391));
    defparam rd_addr_r_0__bdd_4_lut_3009.LUT_INIT = 16'he4aa;
    SB_DFF i50_51 (.Q(\mem_LUT.mem_0_4 ), .C(SLM_CLK_c), .D(n1943));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i149_150 (.Q(\mem_LUT.mem_1_5 ), .C(SLM_CLK_c), .D(n1939));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i152_153 (.Q(\mem_LUT.mem_1_6 ), .C(SLM_CLK_c), .D(n1935));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i53_54 (.Q(\mem_LUT.mem_0_5 ), .C(SLM_CLK_c), .D(n1934));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i155_156 (.Q(\mem_LUT.mem_1_7 ), .C(SLM_CLK_c), .D(n1930));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i59_60 (.Q(\mem_LUT.mem_0_7 ), .C(SLM_CLK_c), .D(n1928));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i56_57 (.Q(\mem_LUT.mem_0_6 ), .C(SLM_CLK_c), .D(n1927));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF rd_fifo_en_prev_r_86 (.Q(rd_fifo_en_prev_r), .C(SLM_CLK_c), .D(n1983));   // src/fifo_quad_word_mod.v(353[29] 363[32])
    SB_LUT4 i757_3_lut (.I0(wr_addr_r[2]), .I1(wr_addr_r[1]), .I2(wr_addr_r[0]), 
            .I3(GND_net), .O(\wr_addr_p1_w[2] ));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam i757_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1_4_lut (.I0(n1), .I1(\wr_addr_p1_w[2] ), .I2(n2_c), .I3(rd_addr_r[2]), 
            .O(n2968));
    defparam i1_4_lut.LUT_INIT = 16'h0208;
    SB_LUT4 n3391_bdd_4_lut (.I0(n3391), .I1(\mem_LUT.mem_1_3 ), .I2(\mem_LUT.mem_0_3 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_402 [3]));
    defparam n3391_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1606_3_lut_4_lut (.I0(n4_c), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_0_0 ), .O(n1959));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i1606_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1574_3_lut_4_lut (.I0(n4_c), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_0_6 ), .O(n1927));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i1574_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1575_3_lut_4_lut (.I0(n4_c), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_0_7 ), .O(n1928));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i1575_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1581_3_lut_4_lut (.I0(n4_c), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_0_5 ), .O(n1934));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i1581_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1590_3_lut_4_lut (.I0(n4_c), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_0_4 ), .O(n1943));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i1590_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1599_3_lut_4_lut (.I0(n4_c), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_0_3 ), .O(n1952));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i1599_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1600_3_lut_4_lut (.I0(n4_c), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_0_2 ), .O(n1953));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i1600_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1602_3_lut_4_lut (.I0(n4_c), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_0_1 ), .O(n1955));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i1602_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1671_3_lut_4_lut (.I0(n4_c), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_2_7 ), .O(n2024));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i1671_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1670_3_lut_4_lut (.I0(n4_c), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_2_6 ), .O(n2023));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i1670_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1669_3_lut_4_lut (.I0(n4_c), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_2_5 ), .O(n2022));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i1669_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1722_1_lut (.I0(reset_all_w), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(RESET_c));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i1722_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1668_3_lut_4_lut (.I0(n4_c), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_2_4 ), .O(n2021));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i1668_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1667_3_lut_4_lut (.I0(n4_c), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_2_3 ), .O(n2020));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i1667_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i8_2_lut_3_lut_4_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(wr_addr_r[1]), .O(n4));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i8_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1666_3_lut_4_lut (.I0(n4_c), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_2_2 ), .O(n2019));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i1666_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1665_3_lut_4_lut (.I0(n4_c), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_2_1 ), .O(n2018));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i1665_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1664_3_lut_4_lut (.I0(n4_c), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_2_0 ), .O(n2017));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i1664_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i4_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(GND_net), .O(n4_c));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i4_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i7_2_lut_3_lut_4_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(wr_addr_r[1]), .O(n2));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i7_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i779_3_lut (.I0(rd_addr_r[2]), .I1(rd_addr_r[1]), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(\rd_addr_p1_w[2] ));   // src/fifo_quad_word_mod.v(71[47:65])
    defparam i779_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i772_rep_9_2_lut (.I0(rd_addr_r[1]), .I1(rd_addr_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n3448));   // src/fifo_quad_word_mod.v(71[47:65])
    defparam i772_rep_9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 rd_addr_r_0__bdd_4_lut (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_2 ), 
            .I2(\mem_LUT.mem_3_2 ), .I3(rd_addr_r[1]), .O(n3433));
    defparam rd_addr_r_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n3433_bdd_4_lut (.I0(n3433), .I1(\mem_LUT.mem_1_2 ), .I2(\mem_LUT.mem_0_2 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_402 [2]));
    defparam n3433_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_3039 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_1 ), 
            .I2(\mem_LUT.mem_3_1 ), .I3(rd_addr_r[1]), .O(n3427));
    defparam rd_addr_r_0__bdd_4_lut_3039.LUT_INIT = 16'he4aa;
    SB_LUT4 n3427_bdd_4_lut (.I0(n3427), .I1(\mem_LUT.mem_1_1 ), .I2(\mem_LUT.mem_0_1 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_402 [1]));
    defparam n3427_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_3034 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_0 ), 
            .I2(\mem_LUT.mem_3_0 ), .I3(rd_addr_r[1]), .O(n3421));
    defparam rd_addr_r_0__bdd_4_lut_3034.LUT_INIT = 16'he4aa;
    SB_LUT4 n3421_bdd_4_lut (.I0(n3421), .I1(\mem_LUT.mem_1_0 ), .I2(\mem_LUT.mem_0_0 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_402 [0]));
    defparam n3421_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_3029 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_7 ), 
            .I2(\mem_LUT.mem_3_7 ), .I3(rd_addr_r[1]), .O(n3415));
    defparam rd_addr_r_0__bdd_4_lut_3029.LUT_INIT = 16'he4aa;
    SB_LUT4 n3415_bdd_4_lut (.I0(n3415), .I1(\mem_LUT.mem_1_7 ), .I2(\mem_LUT.mem_0_7 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_402 [7]));
    defparam n3415_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_en_i_I_0_2_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(GND_net), .I3(GND_net), .O(rd_fifo_en_w));   // src/fifo_quad_word_mod.v(62[29:51])
    defparam rd_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 wr_addr_p1_w_1__I_0_i2_2_lut_3_lut (.I0(wr_addr_r[1]), .I1(wr_addr_r[0]), 
            .I2(rd_addr_r[1]), .I3(GND_net), .O(n2_c));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam wr_addr_p1_w_1__I_0_i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    
endmodule
//
// Verilog Description of module \uart_tx(CLKS_PER_BIT=434) 
//

module \uart_tx(CLKS_PER_BIT=434)  (SLM_CLK_c, UART_TX_c, r_SM_Main, r_Tx_Data, 
            r_Bit_Index, GND_net, n3439, n2013, n2067, n2066, n2065, 
            n2064, n2062, n2061, n2060, \r_SM_Main_2__N_187[0] , n1636, 
            n1819, n1898, \r_SM_Main_2__N_184[1] , VCC_net, n1950, 
            n1949, tx_uart_active_flag, n4) /* synthesis syn_module_defined=1 */ ;
    input SLM_CLK_c;
    output UART_TX_c;
    output [2:0]r_SM_Main;
    output [7:0]r_Tx_Data;
    output [2:0]r_Bit_Index;
    input GND_net;
    input n3439;
    input n2013;
    input n2067;
    input n2066;
    input n2065;
    input n2064;
    input n2062;
    input n2061;
    input n2060;
    input \r_SM_Main_2__N_187[0] ;
    output n1636;
    output n1819;
    output n1898;
    output \r_SM_Main_2__N_184[1] ;
    input VCC_net;
    input n1950;
    input n1949;
    output tx_uart_active_flag;
    output n4;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [9:0]n45;
    
    wire n1;
    wire [9:0]r_Clock_Count;   // src/uart_tx.v(32[16:29])
    
    wire n1919, n3, n1485, n3322, n2933, n3323, n3320, n3319, 
        o_Tx_Serial_N_216, n2934, n3_adj_486;
    wire [2:0]r_Bit_Index_c;   // src/uart_tx.v(33[16:27])
    wire [2:0]n312;
    
    wire n2981, n2550, n2564, n2932, n2931, n2930, n2929, n2937, 
        n2936, n2935, n3385, n1484;
    
    SB_DFFESR r_Clock_Count_586__i2 (.Q(r_Clock_Count[2]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[2]), .R(n1919));   // src/uart_tx.v(116[34:51])
    SB_DFFE o_Tx_Serial_44 (.Q(UART_TX_c), .C(SLM_CLK_c), .E(n1), .D(n3));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(SLM_CLK_c), .D(n1485), 
            .R(r_SM_Main[2]));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Clock_Count_586__i1 (.Q(r_Clock_Count[1]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[1]), .R(n1919));   // src/uart_tx.v(116[34:51])
    SB_LUT4 i2935_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n3322));
    defparam i2935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_586_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[5]), 
            .I3(n2933), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_586_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(SLM_CLK_c), .D(n3439));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i2936_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n3323));
    defparam i2936_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(SLM_CLK_c), .D(n2013));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i2933_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n3320));
    defparam i2933_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(SLM_CLK_c), .D(n2067));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(SLM_CLK_c), .D(n2066));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i2932_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n3319));
    defparam i2932_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(SLM_CLK_c), .D(n2065));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(SLM_CLK_c), .D(n2064));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(SLM_CLK_c), .D(n2062));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(SLM_CLK_c), .D(n2061));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(SLM_CLK_c), .D(n2060));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 r_SM_Main_2__I_0_55_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_216), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // src/uart_tx.v(41[7] 140[14])
    defparam r_SM_Main_2__I_0_55_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_CARRY r_Clock_Count_586_add_4_7 (.CI(n2933), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n2934));
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(SLM_CLK_c), .D(n3_adj_486), 
            .R(r_SM_Main[2]));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i735_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index_c[1]), 
            .I2(r_Bit_Index_c[2]), .I3(GND_net), .O(n312[2]));
    defparam i735_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[1]), .I2(r_Clock_Count[2]), 
            .I3(r_Clock_Count[3]), .O(n2981));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index_c[1]), 
            .I2(r_Bit_Index_c[2]), .I3(GND_net), .O(n2550));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2212_4_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[6]), .I2(n2981), 
            .I3(r_Clock_Count[4]), .O(n2564));
    defparam i2212_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_187[0] ), .O(n1636));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 r_Clock_Count_586_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[4]), 
            .I3(n2932), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_586_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index_c[1]), .C(SLM_CLK_c), .E(n1819), 
            .D(n312[1]), .R(n1898));   // src/uart_tx.v(38[10] 141[8])
    SB_CARRY r_Clock_Count_586_add_4_6 (.CI(n2932), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n2933));
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index_c[2]), .C(SLM_CLK_c), .E(n1819), 
            .D(n312[2]), .R(n1898));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 r_Clock_Count_586_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[3]), 
            .I3(n2931), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_586_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_586_add_4_5 (.CI(n2931), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n2932));
    SB_LUT4 r_Clock_Count_586_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[2]), 
            .I3(n2930), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_586_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_586_add_4_4 (.CI(n2930), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n2931));
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_184[1] ), .O(n1819));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 r_Clock_Count_586_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[1]), 
            .I3(n2929), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_586_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_586_add_4_3 (.CI(n2929), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n2930));
    SB_LUT4 r_Clock_Count_586_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_586_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_586_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n2929));
    SB_DFFESR r_Clock_Count_586__i0 (.Q(r_Clock_Count[0]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[0]), .R(n1919));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_586__i9 (.Q(r_Clock_Count[9]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[9]), .R(n1919));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_586__i8 (.Q(r_Clock_Count[8]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[8]), .R(n1919));   // src/uart_tx.v(116[34:51])
    SB_DFF r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(SLM_CLK_c), .D(n1950));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Clock_Count_586__i7 (.Q(r_Clock_Count[7]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[7]), .R(n1919));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_586__i6 (.Q(r_Clock_Count[6]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[6]), .R(n1919));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_586__i5 (.Q(r_Clock_Count[5]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[5]), .R(n1919));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_586__i4 (.Q(r_Clock_Count[4]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[4]), .R(n1919));   // src/uart_tx.v(116[34:51])
    SB_DFF r_Tx_Active_46 (.Q(tx_uart_active_flag), .C(SLM_CLK_c), .D(n1949));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 r_Clock_Count_586_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[9]), .I3(n2937), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_586_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_586_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n2936), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_586_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2966_4_lut_4_lut (.I0(\r_SM_Main_2__N_184[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_187[0] ), .O(n4));   // src/uart_tx.v(41[7] 140[14])
    defparam i2966_4_lut_4_lut.LUT_INIT = 16'h8380;
    SB_DFFESR r_Clock_Count_586__i3 (.Q(r_Clock_Count[3]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[3]), .R(n1919));   // src/uart_tx.v(116[34:51])
    SB_CARRY r_Clock_Count_586_add_4_10 (.CI(n2936), .I0(GND_net), .I1(r_Clock_Count[8]), 
            .CO(n2937));
    SB_LUT4 i2218_4_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[9]), .I2(n2564), 
            .I3(r_Clock_Count[7]), .O(\r_SM_Main_2__N_184[1] ));
    defparam i2218_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 r_Clock_Count_586_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[7]), 
            .I3(n2935), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_586_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_586_add_4_9 (.CI(n2935), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n2936));
    SB_LUT4 i1257_2_lut_3_lut (.I0(\r_SM_Main_2__N_184[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_486));   // src/uart_tx.v(41[7] 140[14])
    defparam i1257_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i2991_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_184[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n1919));
    defparam i2991_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index_c[1]), .I1(n3319), 
            .I2(n3320), .I3(r_Bit_Index_c[2]), .O(n3385));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 r_Clock_Count_586_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[6]), 
            .I3(n2934), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_586_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_586_add_4_8 (.CI(n2934), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n2935));
    SB_LUT4 i728_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n312[1]));   // src/uart_tx.v(96[36:51])
    defparam i728_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1545_3_lut (.I0(n1819), .I1(n2550), .I2(r_SM_Main[1]), .I3(GND_net), 
            .O(n1898));   // src/uart_tx.v(38[10] 141[8])
    defparam i1545_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1132_4_lut (.I0(\r_SM_Main_2__N_187[0] ), .I1(n2550), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_184[1] ), .O(n1484));   // src/uart_tx.v(41[7] 140[14])
    defparam i1132_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1133_3_lut (.I0(n1484), .I1(\r_SM_Main_2__N_184[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n1485));   // src/uart_tx.v(41[7] 140[14])
    defparam i1133_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 n3385_bdd_4_lut (.I0(n3385), .I1(n3323), .I2(n3322), .I3(r_Bit_Index_c[2]), 
            .O(o_Tx_Serial_N_216));
    defparam n3385_bdd_4_lut.LUT_INIT = 16'haad8;
    
endmodule
